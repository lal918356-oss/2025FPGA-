// `define DEBUG_UDP
module udp_ip_protocol_stack #
(
    parameter               DEVICE            = "EG4",//"PH1","EG4"
    parameter               ARP_REQUEST_NUM   = 3,
    parameter               ARP_REQUEST_DELAY = 27'h0ffffff,    
    parameter               LOCAL_UDP_PORT_NUM= 16'hf000,
    parameter               LOCAL_IP_ADDRESS  = 32'hc0a80a01,
    parameter               LOCAL_MAC_ADDRESS = 48'h0123456789ab
)
(   
    input                   udp_rx_clk,
    input                   udp_tx_clk,
    input                   reset,
    
    input [15:0]            input_local_udp_port_num,
    input                   input_local_udp_port_num_valid,
    
//app2udp signal
    output wire             udp2app_tx_ready,
    output wire             udp2app_tx_ack,
    input                   app_tx_request,
    input                   app_tx_data_valid,
    input [7:0]             app_tx_data,
    input [15:0]            app_tx_data_length,
//udp2app signal    
    output wire             app_rx_data_valid,
    output wire [7:0]       app_rx_data,
    output wire [15:0]      app_rx_data_length,
    output wire [15:0]      app_rx_port_num,
    
    input [15:0]            app_tx_dst_port,
    input [31:0]            ip_tx_dst_address,
    
    input [31:0]            input_local_ip_address,
    input                   input_local_ip_address_valid,
    
//temac signal          
    output wire             temac_rx_ready,
    input  wire             temac_rx_valid,
    input  wire [7:0]       temac_rx_data,
    input  wire             temac_rx_sof,
    input  wire             temac_rx_eof,
    
    input  wire             temac_tx_ready,
    output wire             temac_tx_valid,
    output wire [7:0]       temac_tx_data,
    output wire             temac_tx_sof,
    output wire             temac_tx_eof,
`ifdef DEBUG_UDP
    output wire             udp_debug_out,
`endif
    output wire             ip_rx_error,
    output wire             arp_request_no_reply_error
);
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
bYWfmef+IesTiD2TYYSL47unPhAW5jIZCesukRoHVm14bJraRuZi5lOUH6KbI6vN
K8Wd5hWhE9wzLKt98ZOftrwOIxHppC1bvqv2lWKKjydhPxEzKOIeOmHeBkwvcsd+
5/b16pq4lG533NWBY/wR2+D2L84bEvTXI/KJpyhU3UU=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
X2QwGnjpx4j4B1zDmHTZHkhLsPLgTFVPC0yum4z3Xei+i9CkVm0pk7hP1xTzNQlA
Tmc7trkZx2U/0uqxDeJShxMzg3ClIuxJyIm9g35g0graw62qx48VaRpNFqeIsMy2
Mq10W3Lhmo9Zl18t0god0Gk4x9eq3OfbyWbB4ovWE7A=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
AXH/IYY3Nk6K9QPm6vKBoDuYlD5DLeHEo1in4UBKj2fSdGKUK9mgq3W81evlOfXY
YwXIVSVDiEtJLTY5LQz2IdjsPUiERnA/W/tnMc+ENpEjvsJOJsKMBd4y4QkOQmMi
QZ/4ae4nQc/fFuxOJ/ih5+DJZqTsyGbZr02K9rvrdSm/tkT7XVLXF2njqAZJr3w2
28FRtNrFrpiKEwANrj0QhevX3ZECcjDxDQBAay9M5MPOkd2HGdu+3AVBlefnGe/h
zddSi4cFRij6ftHC770ncZ9Zrb64YOQU5oZgPu/SqASxwvtAR28sBJf58ITGU4BV
HzazXWkSUM5NDB/jWy8iQQ==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
RJ7tqQTOTbhVV7pSbA5EtGh9jdjFwD6/53Z6qY6259C/e0a19VLk9EvE5x64X91o
laYq/2tRvV47wX2KfGqxAWhMnLFRSg2HeB7BwsIgdG2psLvOfdTfn1r5Lwnyj1Zc
1wy9LMZYfNVsFhP93xnB4X1vRR1YgCSducMblvcVZ54=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 15520)
`pragma protect data_block
TOXCjTraDv4cLYzZILt67bS4ZsGQCXzWl4tWxQO78iuhA1fFbGAEluKvpLZzLD3m
XX/qEKMddrD5E9cGC0SzCkLqEX0zNm1Uwx4v3rNXVBlBziD+PbEYhfsyr3byEg+X
u5r7ba2yJs24l8IW8Fm0hUrGyNMZtLy4PxuJ5xDk7no7khpLeD2bNMj+mw52HXBH
R3MUUAJfkQOgDrcB1BOD5k8pm8BLsHeVCIMjolOiI867blUm3a1g5LXiHu3oPqrw
ThK7+xF9F5RuYEHX474Z7WuO1zqZOf/AsjQeSISqcHwaScvFnxQhbc+WH8ElLCWe
5NgB2OH0t/H5MGjrH65vdaQBYHR1F92BGuod2QaXRL8KUMUJMtWN5w/zAfaOC5N3
nM9m1+5ydnuq0KvyojPfEqZbHGN8ojYvxQ4CeNeruVyCeaNqYkBiZEyBGIEHPZ/+
KionRr8XOn12YgvEsrVW4zHC+G6YWs1Uau/k3INRy8qxb2+BdL2f+/Prbq5L/5fY
bn9USgVtV6MxWPi7LP6SgJuKeAAP1+ZSx4DaMWTRHz7naOjxgQ0n/lSL3i5Yg0l8
PEV1jrTYoAmg1WFhmcZfYZzTk3dnrA+3B3b1wlPDIC+FQqR8Oc9MvJw0xsdf0xwr
C4+sNMTuOJS2gYzRwtEned+4mZo/gvldWet6TtefRuzZn98i2pa+KKaLj0wSEViJ
01pp770Easxum/UgeD6H1r51M+ZVRVjVT7UzCr0Emf4/NwqwyyxKJqamb2eNpzPy
HY53HJyfg2dk1L0I4cHW+bwdvo/ffqAyJNaSkCu6Iy5DHQZyu6RKRf88fZ2zAO9n
ZKs8Vc7SRXyasZb9NpWvX/lwyK6l/dgxu17bTZiVsp16s4DOxsQenDYPNHKARg72
bFWylE0lh/hKoU3VfGsE3p9MO0nw06K1b/sqDuMzrnqtrXeHvueJGxN52gzzFthv
YQnO9jxDVw6BTag0oESwS+8Qk8RMYLLslINPV4Mspc/8ldQHk4sb0dyg93+EkmUI
EI6jqgj1wzjPFpDKqEeMi/nM53uzSm24b7XWHE5G4Cg7FhD1/XfMJ31juZTCa4N/
TcHmGyL5WQCXdoLZnRKjsSKphtGDPTzWnL5FhJ4WtubklHpJF+iH6XzGl8FUF1mW
PMeOpgVgOcjkfEju13ElfeuxWmiEuWX7sYg8HeVbyxKcDnZUNl/m5Xi3yJIFh5fY
vBS4iXrEdXloTINTqV55MNYIf61GOl+5wI7AqOIRflCQJNW911NKH/7ZNCy41928
yN+nXU50Ebci0AGe3wJnqM8aJqfakcGc23D+XcnXyT0PTUofKEYpQSpYc1E0kJj8
pkwLf4WE3BUd72kfN5c/pwImRxQeTJz2u+UQUYhRXEFIJ2V55Byc/HYdbe6/ZnPF
MGQqukjF+g5GXOey6Hnn0Z0gvGzDYL9tvAzs71DKflhd5Fm6ruGhS1BhnQuuXU/r
Rn6/jdvhD6tSWIYCvu9DXN9KLFEf/+fhZx7oIFZYqgIxOLY5mn9Kb/SKbOoMNv8W
Cqe69j63+x0SSV+1TUWOrADUmFNmZk5rNgNTXXfClcxC5hPdABN8PX9FkhjbDd4r
LbH0rDHDHycJwXsga91tpZ2Ll+QjmC84/Tk5vBW58CjNmtTDbqp4033wHcnOY4oL
nJcBclpdtXMwjFI3kRGTK6mJ5KqisrVUCW9CHSVZGZrOb+vI1KVhlnBAadW45X8W
VjVQULkqmaVLHWcPCcsMDJOBwiidGXDMhEiOc1gJFOf1V+Xq26z0iA1yDMRfOR2g
HckkWFkNvImteOUg0A68M2YTRxprHuzqU6lxZ9G2Di5iyDUo8PQqC4Xnf1Z6E/3a
DrWymuWbnnnDf7OcCdgjV+2lXb9LmakCwB1K07Q2U4mFq2GLwThAnjBD3QprN4iR
mGElFCZKtF5daHQTBJtSbAyKM8nj+LMlJl2wvn5+k2Co6FV6ybN2a5ZBuouNlgKG
6apcsZGVvRDdgH9Rz3bcLyJuHK6IiyOWq7Y0jSiVVa6Iaoltx7Pppp/kpIX1i9Yw
CgeVetJRb0DtL+8qfC2giouKXib2Dl8ATd+BL9orL1+4X8uidE865U/FA2uHg7Jn
qDKu6KVDeCa3IYsG0N8Ac8tjODFE3FmIZNxpF3WvQBn/x0lgIm2LBv+EPgRoa1fs
xjIavuUecyy0+47uLkphOWew4ZXV24giQoR26OtXaGn1NZ1SNBlcHLtTOv4Vhxv1
9IAI6gnLoXkYqJxjtWssV/HqmpVVSufEaa3fqhamAuUY44GrCTYnOqIudPIl4tfb
0fCj5sCo1cxSQW2zOMUvlLBOEIfXa637JJa6WvoUksR9j4phkzNoyYUCHhUwhGqH
kRgaf1jIkXIdRuAnyDuMbOOwM/3ensWMAgrXW1VTIFFDYNZbs+ZsamCIX4h7MXCl
SZfjOZfP8y0KCArf8GHHsR1G50n2bhFo592VEF6YuPtzUOpJ7KfZzsaQvtbPGrDF
Jn2uiSxUBmANKwRVI4VwSfuSWsAe5eMZ+R+hXlFrlXXPH9ppgy7BaHPrPZX1et9D
82eJRpeI4mGN9jJ8QESxv4tluaNtYGau+4ZsTebeecJ1B5oVkNexq7xQsRzm8LuU
4rFnci34vGZRVHK4n2M7OZQedvoLQrrozy93GOkCqstjKUrfzDQzLekBW4cAw5nK
EpZVBIxtYVHYCTk8NoBES90HTVcVww6AvW1pStIWJzmOeQgwf6TpBdsW0YYTUd5A
nhx67Z0zv/hZAl7NUI9kPXeSr8t9HtJ2yV9+iFrRUyPGL7w8gI9D9zUmQyAJ2/Kt
jr9qkc4lnw4/eF+2nDU90ekNVop7coLWw38ap4PrWQGiI5utdqlnzTZZo9g5NasJ
ExEHGuFJGTAKw8n6OtqPeDwrrEuRvP0T4xqfZ9rGrRyycDQ/yTJQiWmA3TlqxOQn
9Q9I5XPA7JYbTh9ffzp0LtDswiGi+BMdOit34rCShqSXbSCviaDTzBi/aJIgoSHn
LDgDuHCelVZgcmigTxnpiE2B/iQZHWgdzHMik54Kfs6i+ydqf3Bg3bP2aOOGEo7p
mEOXr9rrU08v+/rezbIzj4FIG9rLJuBJ/NRkYYYEip3JpxdwMFJCXC1Z2Ybje34v
OC8NAUq5QQyYK2ptTa7QJaIxkbAGS6731/rfzZabYqp2LJzxY5NkXiPvhZNBypD2
SgvYLJ+jdUqA4GuHXvrIDCUUIrNaR22qCNBSOdIl1/SrabLQbh+L1nzK6HAPN8T5
qFMOnnhPLlQSe+1kHIPB2jHl2Cz5cbrKK7wqydDQOTZkEADal4YC0bPmk9Ybghe5
zrw4DoBJl0azzv9aVCUvcKFgVyEZf3ywNywbU9Xfy282wXqSDtCkOHqVFqyKinpg
ndZCc7pk0tI2jOSgcOYq0DNFlJ8GRPbbK98kAvkTEuY4aoGcVMXSCvgNZAW/EpGj
ptfhLk8pRenZoRjop13K8/WDD4Km+4tFFFfAYc62MntIFprYGs1bsQx9Fi5m54rx
vOSmXMJhv/Z8+rbf4RzD5QrLRxtbf5T+5VHbkrEwNbugc3Ex7i+qccoXkqp6EaZx
FtO9f0jwoYcofsJwJtewuTOhsMZiL3E9dh8lw3yKyV9bA2BJrJXY8dbCJNL881W1
QmA0lQPrne+QeHpJ00wGxKYG/voD7ElzMdCaTYTUX686vVbs3lCSdZpeEX8ugCUr
BK6mXFNhNPgSBEdO3eo4o+vRrmnKtjSdEsfPru2ZUSFNzI5c1HB442UlEUkTshTQ
vFKZN3dS4LJYS7Apy/9CxnVhdHB0IX0+h5MPM+1lwyXn+odZ9Sleev0BePhk2oXJ
Tsvk9VnduG8XMPFZmWIUWWwbZeFm/qQPKLKeJmQlgybZtuFeEAinvY9+54xWwpdM
ogWgPZAjzc/eVBhU//M71nxHnNQ9ycEElLhV+uyAPE10RLztIXlWyYtyjZcck1+X
xPaXUawZ+5Qp2J6b1faFCMrDN+2vgZL4/mL/NA0bAV74v3qC5VHTCP9iwvHBLEzD
9QJcQK/Vi8Zb1xt+La4ty3AXO5zGU2N0+OybOvhdN1c0BSRlZG5n8Crobo0tFMzW
isW7Y9BqqYrOUknS9M+8RQhExBsJEYwj7NTEZi36fXhd94U1lMFtYJ6j41EvtglF
TvIER1Rw8LsoPXzZHSJ6s8rcZK9Yz8xa4R4T4KwsWAHPyVpcfgJ0copIj+iE2nqT
gyW787sWN1uyg8ypeemnf/YMTmtfCX4ILmyzZv8jGQLDUTfM02bACRV6iuEF15yJ
txhPHiq/4QLzaCfWNsiNSFKdgNNgMog3+vdD6brffv4ui58wgPSJNk52ohsMsBlr
5XBdRrZ1fA69FRXf3jruXvHRFmD9Cte87I/nR0o9nQvGdW4+H3EQIypiGQsSUKqZ
0s0S+smapEH82DMtrFr3TU5Z+zTWrfsQqmp0yGOM1PK55Os19z1MqZOqlUpN/sAw
jpqsI1a/eWzqHdvs6yeXTOKMEviz1aJ/UBTiAicF/dhKvC+CMbYJpTF1fZpsscY1
4iaCSuz2z9yeAnL0DQR/81pe/+VTOqTy26biCWuZiH5WPpqGT6OA5hDamHHMyvmb
XCDFaWmPwg9eyBcfZiA05scfh4UPOrfPRuUAu3+T7bv/gu0udqobX3klKnpoXG5F
cg/bFcVyldp8Kl88jnifsnggpY6ZmUcGTMDcMnlag7/RXwFis8OIW/7bH9d0zkYN
oo205tDLp2VfXlzv3tz7EPypCmCAaba0yHtNc7SJbiN9eOto8MkWZuwW9F1Xhvyz
2nl94Wn261Cymsvf2s4CZowpBktRKG08DW1DVwGlRyK27SgE9bo5OV7ITViwCVff
dXZURI284iUkVLoMBl4SfYI8tWyKCqEp3CarzTcwDtXdrbzoRAYur7BV3Wn94WX3
MhcZP7/2BE8AEmcmN7NGWWGGLz+RJUJZR7v7/lBI4ds4GEXY8q5Qrp47PJRoU/VA
oqYg3yiV+7SIZq0EJUXM75j+E+0xjfKlduYcGdokZ9xhYy7u1k3P1xYgamB1hqVt
W3vH63Su2sxVA7deAQ/+KhUe4y9+FIENuVPQjju/bxUiz2N8BXDvzrLvlVgE6OWs
kR0UVPv8LsAMlErR23y0MFjaWFdyxBTjI6dcBcdlJAgDubi2WOHzq9AWHIduaVuN
mTx6FCmhjV6uC4IwtAK23+XuY4P7hQj+YbzgizevzAHaHIstwCvnm0O2uEQpPwHW
f3J3jDnAEG2IUwO97Q3hVOp1lKjfYZvTarwh9qsyoN/xAHwyJx8x3FqnsfYLH3fL
W3tiOzbfon8gJbyIv3NNxmm3t/tFpMS9FD8B8v5twHfDD9f98qFBWwQHv4W8yv+x
evca3LL1tp+9ndJnhUVlut/arQG/Y4xy7LJnfSDcmOk/FucDSREmCYemSYWLnUqI
ECx2h5vmjUL3k7dP0DuJf+4yZaiQJ6wdADlG6+hMb6xZiugUR9H8FisiFTL8hrKD
1TacNG4rekShSjB7uyLFVzNG1VblILjJt/fFEtqg3Rm5cWdAfG3jnlUI30OUBXQu
wimug9dHp+biHMz7Fm1XVp/fnzjmW7aKB6DW2HFbjzop35Ih/Acwm/F8MWEWM1Ni
Ho9SXO6wZNrJN3ebhqaxWtZECLVhL2stNkG1W/HA61irg9vOmOVizpRQx5hmKbkU
r/6rUPH0C2pl5IAEmVS55ipgZFW0Wc4Y1U8ObMlYjZR1LvBYto+aa6kTpaswlNSY
9mpJDpMbYx9ZXsvEXyUjZhm5gvrcU2hwYZQzv1uYnOZ2GVVX8sXffNQzNK8GW2sl
GVMgio1A2pPG9JaU23zaViwgqZjWSk9j7wG2O9aP/dwx/DGLUZpI0jem8VRaiXSZ
2hD4YoU/3Tnlk/5uZsqBamYB/l09t9JAt9P2Z0Z7BbzrpMwllQkaZL6G88Eovz0G
9rKpt9d3aZ5jWnH7bfP4tVhTtK6SdLLXqHFySHuTWLMC43tB4d+hQ/7Kg+09iMDW
WSO0OxPpDW3U4XWz+mXuHhYPFFchYaYPSc/CQhDq8qrOdYOgoNKkcwLBtgsQnmSO
LrWG/Ft4gm9WF2CUvlfoVoRrZW4zUzPlVNeEvXo0MWQgFOty+RKZJfPDHJCtJQ5h
jfXP1D2V6gNbYdccBpGpg5BxmV6nV23m5+b8RjY7Q/w7b6gfvDhgTstRmrlUWW0F
nqXoHTpzT5s46x172oe771Zx8ZYedmGYLg0rzi0EV9vCaG7lMbMqIZmY/Ao5nArd
zJPujQiORGaW9InVkhi/LhbSQhoYDp+KA0xCLUp6qa8IrsM6CI91qLmOWv+mNIDY
dhozyXS4QeORkvkFInwdiiCMDGMYta012+eYK2txm5RpNdlY7k3NoYyFRd96xM0B
iBumXvj+/krv6F1K+uzHCTWta6RetJXCdsmFyJ5ffgd+IvPI8LX7DhWK/Vhx7Xii
wxEl+1fdP3U6xMd/V8FqfvCQW+1MgZ9AQVbuAIneRcq+YhmDFh5Vebj4T784vcjN
h9AoIQ/OHrsmVg1lqrxA/W8NpdcPd1d0TPW13uIohkOy2Yf54cKUBK+lbD8PPt8A
KlaE6AySaYnjsmYE1fScFguZ5xDzLprJpJPKDAjjRebQu4k3UKaq/VRRwdUFlqAg
YgiN3a8kd0UVhtHDMoDWhDLF1aDA4s7iCsFg1Ve0gGyfLYolwAttjQqUekSGHA9U
LNY3mWzBp6S2NJZ5M62daMVVGosQalgALU53+l5heLUREcbjY67achhn4HfQSU+F
gqk8icdpNNE8VbFOu5/P/60F6dCT9DGxPoTIcwxDi8al2ebLPxDPiJnFjXJsZQRg
KCkyPtjqvk0ev2lpV6hf1LjS/Q139Wp1mrotQYqE5lJpL8a4X1+Hq6NYGc/tRICE
1xO5OsZdb10Ip67C/UYFzAW+vTxS8rfmVUXE32D/TPKIyKT8uhK5nr6UfCN7zV93
FffmWGae0qndKra2D1EtVsy1PktVzi4ZoNxabmt0LmZq5F/UIFHPcLkNAw2uYIC+
2TG20A+ODuyOzTEu5POX9MQTfpuDVMLUsubS1fSYtT8BDcPflbzp1Ekt/Nn6Mw8W
Oxy3qTd1b2j2cm5xompSbo0Gs2X3ArcYEXqTmv+PalM/S2i/7YG19sciTiLs2lId
H13pb0u9O9+C2bIqd/sE59A2bhVuitPYWyifzT73PZFmdQ+tcdmLTZdhr3t/mChp
qOAKily4vmcQolvUuOi2g7Leupyl4pHKsZrgtVsgOZirwVpS8Qmi5dDaFh1looMS
rrsQVxWJNEXL6A8OmhNVPwTOcThMZ4Feh0Uwf4Z/yBcV7XsoIgWvtDOwfenr4TSZ
HC/TYaJchJwqI8gp4LA7YX8mmUc4lgcH0j1rxjUcihQKEBOQRxlQTU6ZdOAd5A+x
k0TaoJ/mPNCHFcQynKtTo/LJ6uamcWKbmfiibcOgS9e1+1S6Qqg5iXPn/gYpeRna
32DAlB0QScnsFLs/KjVyuIcHSO6kAv9zk/Xp5fvf6jHZFnzc4oMvVnT76De2NoaF
n0B/46OPJRQ38XoDsITQj8ASc/xZqjv4m3P1GU7srquHafCca1fNKazfOvARpN7B
lPZ9tegjoTpE5wWP38uB98cSFfN1B6cj/MIAU8uM0LvyImmnTnJ8U9aq8h/83nMd
5U3ZtbwokY6cjwmzEN2F2zj5OeIYmDpdkRrx0ekBe8ezF84PjTwG4JYiYnCrr6LT
QvPpm0DtcfAFHzJJblp5E+0P7533R6t5ancG3XLwq86tcZKg8/bCP0c9nyN97+MJ
W4dAHPGth6o1dQVtJQ0iXYhWRlH5BhXvmOFfv+Sfcb6E1jaUgwz9bq+wc7vI7GDq
vk0whZpk7LHWTDT3tDQMC4R9arAuhwOkQrqBpPmlr0D8dkZvOteN3DrKo5NkdHT+
Gw4DJqIjn4rNAWR9IsVMYtvJAu75s+JZUe9yR57g2Oe6MSvzpq4XgJ4tprixQGQ9
7aZfhjviaVv99+CBylY6iPq1Lu2pAkMUfrYvQmAqXG09RG1IoN6DF06HUXJs0OFL
g96i6tnrNgyWHXcDFYrRqwcRv+R49MGKNEq/nobJa4Te3EKU86etY4JP05JVwj0p
Vfi7Vk+vECkZOVP922OGw0Qsy+Bz6z6rDvfG1Qj2UW6RXRahb/pn2/r1ZBsVIsh1
pKGv33ou9izzXqsNJjCnw9qqMEfBvpJSBoVqt6X11m0ADo+Lrt5sUOQb1ZFaImKk
lp5YPS1Eb31EpDZht/hjyg6EnxWyjhzFo8RlfX0LfszEARh6c1bBm9bvdgKqGfLT
s1HIVH1mpRn2n8XOCD8h+PEvXDZnhUmBIiFq47fraAwEqk7i4qPgEhvT9scRd9Sa
xVyhsGuPx9l454EdGGJqP1U1xQEJyH62sldPA+Lf8Nu7F2FewDMUp02Qa4uESMCi
KFwK6FCVgCMlnY6+etC+yPT+KQLFgUAI3WTecIrNXw+l0pKvONDbvXtlhdfvjP+L
qWDsmFnGn1+Ttiwz73uxyzwqzh+yZJkRNn4wiIIN2lQQMYSa1+Aif3ogzvtOjAid
IDC6n/YzdS3d9rNeHEQjaBrD6pXKJw6VfuX7IlPNdgx/NQWtmpuu0YhOHll0JnPX
dU56hmt0dxAX6adEv1uIC+s26g4n/IZwMegZ4KzUtTR8RUltm4LJY9JqucD9BGhy
XdcBJhtnnv2Bt4OLMPgBQt6Z9N/6r7iYey7CytWROgMz9RPqOmIvL3OFWawakOY/
LjgP5fOYtD+RjvV3gpZn3bGqRNn0qa+3tG9GZSgD5dz2y2BHMAcdmgBtZybttU4O
2POwWkl1zNZRNLnSazDhBxfw7U37nIlIe/HeqJZEo0JFxkdAS710KLoTGWwEl+yb
Ux6epmcg0MHIfLboxXqcDNc1iwLklffCN3bCOBjRM+SBzioGqu8nU8kXkkVIKS04
Qu0g0P5qOUkWH3k42UdFktOdyqINcSSo9ERicd8Gd5u3sm3vmvvVPeceQtxIDAeu
PUBTzG2dDY07ACRib15BXRyD+KTsAYyeZ2ZRor8Ad8fDueVhxG9gs4/dCeuOW1LB
I9StopbQqxaV6P13m9FcR5BrPgxuvQzv3LiyHvBF2IeTlthZvSxEJpK2/bwdLhq7
4Tyh5efrBkBn7QUfzmQOUCqkcljHjbaOFoe4uK8DjiywbMsMh2IHSUgRioyH8TOX
3PDB8bxdLlMK1V87FcSPC5RKEjXyHOrAIpJNRcxhrOWmXCvmyLWsXGsYLbJ44qch
MFEPys/vMzBpy5exD+rZpp6HAtHbw1aAOSbnrrsECoq9P8kuIsvHmK9eufgsAliv
4qEr2RAIY0JZhMpiZfxtlz5S7NKPKFvbSnhDtVNe/cLXvOg5ZRP8Trmo3EdqH0Vt
od0t6YEkyeTdM6BrWXn+PHmyqk6jDQsPrwrGGYTFq6HpJD5iIioJgcOgd1WyX7o4
kWxDcfstr8m0XlWzauoLGrJYhRYq2UtBcFNd4CTJv2amXegNoz2KKcGb1S4Wwytt
sH+snRt0dYIVKEUU2TzdBisViWNMpub50NNgIFVJJ8yRDuiiM3EcLox/xQ8CYS2k
t7ir0ttY6HnqP5R/Zwon67wsnm2d2USrEQRqVoyJnJAAnz/yZpGnQ42y4Udosu3s
uI9080oTFWqmupDM/7gde3d3Do+C0A8nMYLNy2jj+KGMm13cXt88NDPdlKlC+jXK
S7MTj19Ok2VfjKVlFPLqu1S1yoEFZXccBHH4EuGV4UvMAUH9qkJ9Su3dnlrgifVo
wAo3ldpa2vrkDNKAaGxTtr+R8T+w4WjpqGu7axbj911y0t1k/2ou2P1XgXnGIeFy
+44wcnZP6QA4rGEeaCwHJzQVABxZ5oMCkq/eOB5XRpFtO8gfo1NAKrmcHWeZ85cf
rwBA/VwgqWaqoO3+Tx0KpaQarjb6aPIlIwVVJVb18lhHWIBtiADY8O8S+z2xXt2L
YYy5HzNIog5RIDChUQGVIhli2jwAUmelOqOvZmssp8tq3TrWgogUhL14tf0brLKq
aiYTtXneqhMs580n1TkzcdcBhEimVBZm03m0Kas72jy+4CtaDLyfLvU6pKrWr1hb
dDTP7MxrhUmySbR2IN/irzjV1l74mJA0cc4yAYXgQUsp+1GSK7bzX/p9fjx2KaVN
80GD4Tt7KKE+A3SCizPyFPVsZpRaceUGNkghff7IOCkpiEBO1XShNuS8CkSzEWK5
f2vlCuUAuM/zGNecA678aRqFRqNAEn9lcv3kTRf6L5137guv4k7Wl4JMAW3gIz6k
u19p+ICFvm85nTmlLnnPOYukAm6nI8+a8DyOAWcuGelQSEQZ57Lwe8Vuhw2WpIXC
j9NIW1Aczdw96Jfs0+xu+qEuKEly1fDeTBllA0ShK+mheRd6vRkrCA3gAPdq9XmG
O2uYMbDGmW4LCZ1CExcbzpiW4EsF6+GLkYCtobIVQv5qYi2bpFq+CaMzusO7muHt
KtlpBccyGcasA+p8FZELxsy/0pRXNpMmC/Tpx6piVEJxl5oJzSVscTQTpBaBrAEC
9BxrD0qSpa5CAasWOxZ/8qKaZu91px4NJsbbMruc/+7PW5+UWKtcGtua9BDnCER8
+0Gjd6Y1ATqZmaF0Fn0q12PA2XCRyCY1cNSLE9nZ3hcaqwr0JPgZCgWEEnn4AtdP
STs4sXmUnzuTWP+wozdA0xeCCtjK+QB1RrsrkMABYKQkdKVYcpkipyAQDat7f91J
ss9lxKcGvznwyr4ccoakWZXOI+Wu0ugRAvuME+Chmh5+SzWrsoEMbiWLbHKN7TVB
h8HOTD6i6kKgibObTMIJ9611XI0Uop5j0vK6g5gtiFld7bCD9QBKH21wqJY6g2J0
adMfi/4hgwsa602lrb6UHvwOp9WxOeiMKh3zg/87Z8uepCS9n18JtfX47sBLGaVK
rLl01NixI4DC3wFw48uNXkNXbc4OrIjS37qrBVCbg7+W2j8dHrbCmxQ42g+mRvlw
AVbvglaIunUnpHAoiucjz5gxZSephOQvRE3hh8QuDLBv2iCYbw3HhX1zs9poLqxk
YmHrIcZ9l4aH//UskcjubDqtTZ4/x/7+nDo/nEJfxs5Hs9nGOnUD50ZdA+Il0ELi
uZSCQPVmtN8yQ0CTmeWTDsjIIUWzYpVhIwRSSUFPrhJPNe1Bw8OS5bAba8KGVEhC
CYdWL3AHp3bK1DaPgcR3P/mCwmlNUOBv///H2HNTJbtJPDjyH1FPAUEzdR3VU/ca
+TBxoMyv0QeY6ltJ1/1DnBssuU+h/NWkaCQ31D42T+TbujEMdf0rYJYuWNxqkm+A
EKqMsjPRTxYW5gDxLThcUFYKhWahcAf5wQzL1UPo1rwL9ST7mDCy9fBULOjxgq8H
ZZLvJyExbnlOKbCbLvXQ5wJACCo6sPOC7LPZtw/X1aOEzP4FObssHOCLkUg3lT+L
w6NuoB65vPeTV/FkizatEDukfrDuBkwWlcZGTy4FfdULbKvzjkaYwTg0ZAAVUx2N
L0AX5tF33ENcdy9bXk5pvhDpQLQ8LUki7oEWzokaVcSzZcJeUnHrJ84eP1e+ipUD
5ItUM0QkoM2+1GKbZBC6FJiCp1JVvc6bC1XZfxQ+x06OZ2+SeGEA3SfwIne7zXb3
Pj68fAvIFGeMVkYz29Au4DFaucPiD5Z61x9WvgsXuNATp2y5NivvcbGOABno1qE9
d9sM88ktNeXCSmt3Etu2sGM+eXYc5NCfHtx7OBvPtByBNISGsx4lliWH13Kg0vod
q7/5HYLHMAU94uEWCkfqtiK2onurn0pzKKezwwMYbqx6k20bCG1A3siQBpOfpeHm
lPt81tNZlXtY+x00nKI2VYvY+JpAz+gVefcPky6L3jYxLJbe2uTAj8SJs8SzzyD1
NWv/u067J9WQMLNkqnUCVl0g9aiKinnzWtokmglwEEFaAKwsAIX7TMTxydjpATeZ
wkNOVl4BmRNExgjf6mhj2Ja4GOPKaHiwYwyatFzgUKoHQHI2MXjaoSIhc6eQtVfy
u6+OejRNH9Hg2I++zXCTE5FL96W4tke5eHGmyaVmQ+jvedj2hDhAl32mg99wMjTJ
MkyqfbltSyJJOVKrWiSeOn3DlClQUCEY4oH+VIc7FK/61W7/iwrhbwcu+vy6Ek6m
xym0wMwcjCeUygzQoX2GFV/VjetIwXSLKHt2XBjJFAqNB2sTdRHXAQDdbJeiaLF/
UXMVzAGvjos439O1kYJqowjVYVYimNyMPSKPISDjHeeTCTLmDzCljn+90wHKdNdI
JhrwcJ3N7SqUP88Tcwa69S/thbnhM7zL2OgypQ9wqOudO3IcbqxfqUcd5gd+0fkL
2tQf0Qg84WXqqwnTZVxS3vdbXk93iWcnsokLf9OJE9MFxTfkpFyvTd9dYfMRVLcA
Es++6F/9W0bCpQDhxVP/gAUATWvZCD8NsmIj10hSUASKiDm4usDpTLCu0FSoeVIx
nyUfMvXfyW+nDj9qDyHU5BIqH4BusZU2A7DJULUDhFW0NT9hz/sxNsFDZfS5Rxbb
f2JsUWogbYuVV88Zm56Fp9QJ/iPm24DC7IaBOO69+KUlApX09yNeC7OADajSBfWZ
M6WF+aTFP55pm81lDsfaZbm8dEhzqGOlNH3fVBQzVfTrXzD/yz1PW8qQ7z0EOIcn
HDq98mcxMVROP7IuDKxGSiuSDzH1sNt39dK3+vBWSW5WIyeODDXPh+tGQBAZ4LDs
IKF0y+CJ5siBrJoV9RIGbP1plFW5Jkm3iDNVNpWVD4hAoyomEmLveE7KCJx8xnAh
vKVZNwKsBlt8O1JYqfM1NdAjCpXec6+7uVpMX3OTRKq6/Hf38qH1tUC7si37zWeV
1GHZeoLwP3mYus7xdnIW7o+huBMHCPLB6MB/j8/Wc6BQaxFIuQXo+5IBXbGjOMe6
VU8eR4IcSAZ3gHmlYxoA3GFb83FcAEvuc56M00PN33pCenc8QLXqSNrHOVX79SeK
zMTJOSicUCwDbCtYWw6kFcWC2bO/oXtBmgNtPrk3F/izuxheKrYSKwevK0PFNdFx
3w332a3OuMdCgDw7kEDQE0ksYkcMG2VB0uFqtCtKnw2L6lN6aZvKTW2sb00IcjgW
pO1/hbgyyxJvudvugei54fnc3582IO6YxEN/lvTbgwHsAkDk+wRIigc/1h9rxqvo
/VGj/xXTluvIDaZgKqMNPn3uuR3SE9XmKE5DhSeGn2HYGktAAykSo2t9eJspy4Vg
cLVGCiYL9ki0FPWo2IdRkhtWsdwwcD/DN4hoBq+VAOywuZafeLeqPP/SxlMDUc3g
afT+ClliauekBECQzbqmvoIEHUd8u02dMwJKhopmesgwSPeNNa9sP4e8IZqC9IcW
w4vN299VJQMAvI4OCS94yYQT0RdYDxjSkljmTbKWemu/2ea7CIdL8OJQwazZtMqY
Df2P8Nhke0yiLHypFueLSTo0TcWD8UK6QTuUgqsUZJNV7fIuJ3uFqMEo/AC+88yH
SFODrmDesXCLRni+TnBL8kk0JUiEeG8SsMkR82ThowYRCQv9Ul2el84Yu1egOsON
p3EUu4kYOPUsXzMqNAoMlJUjhH9KQvd1EEk+6aGoedI/tVI6oSweLKOLHJ3FgbS/
ozCeSuM0G6lX7meAg/iogb/zloc9msPqDR+x55A96nVHzXDAx4Tmkvq8NNgbjF4A
yvTgKlkoWFdJjnkYhRJgXgVuBmgRsqZ+FsHRe5ge/S1dMUbjsDtlTGN3VhvD+4vB
yOkNOm4iavMOroI7PaeuBG3xCgWWa8EmywtOXeZgcs0Lx+igr7PgOOM9JYPRnnSr
4ye0GUbqAtTE+8fpoofeGxhyarftOOK5k/H3SuGh6rN+BBFU/W4lNHeyEckNEi4Z
+PmnTp+0V8JPVnVSdmK/WXNtWYprN+H1EJpc7Rh4b3R9TEXucpM880DLPXSbwLsW
lcvhCXohBx0k9Q1laNDxGiJ1YwC0TZw4h2qEATF6/lPIpMUUPR98q5FaUk7/ZdSh
uHLEpORGYmRnap0QNx1XqXw3f2ZhbOANg9dmSRuKVZYXHf1JqjaEw50Yi8qdWpT9
aflo4l6rncS5QmJjxsA2Br2U3P/mpnZN5jCOwzU2H9pytz5FXT/T5Zt9e2txsGMf
KEE7CoNSlgkVyC5cYDOQi9JXV+MmniLqrWCpzxQP6cec/SPmxEp5etMUutg32gWd
0IxN7PnM0fJgVqYnNsrJ8eGbhBStM1N0IAFtNBORfeL7powQ97UWdOq+R2dfRArm
MLP7ECcO7zwQ1w6qzGUpJmXCoZvjMdC7PiI7HORi6to/0BxR+GfpvODSE3mGc0y8
dyi0ndBntxY/UEtQu8PwPaD1uWGVplCt3k49bQXaiWsimvEuAeJc/7mTt1QWcZ4F
jwXdKsTPVxi8yfcPnN0GYmTMQw4iVpE30zO3y3FlWh5GhnqCojIDkaIn+hrj4w0E
EYwyJdpVmMDuxqBkva9ZrGB+mLufTppyMg7hRyP3aMqImeEVRaP72EUZk4p32+Im
gj4YsaMkE+nLdQ5GB+M4Vp5+41JTTlQ6j5+DhI4W+5KcncXLq5+cikturKcuZ5i4
6Q+bQxpBCqfd60QIjHDB93k4B+gm+FPvc+0xwO09zDRuP42bX8oAY7+LRuqG7XS5
W12OAnxBy8hFEMODHHtX/ngMGj1WrmDMqaVN7uzEbHgMEgqGAYOLHNfc8zDBCFCB
8wMa+W9VBmK3T1ISH3lmDi+9u+CPlhPK/hfQCYCjd5Gkr0XSatryES47RGUihXAk
XDAJsJgBefdF6EGyYxFVLWFvWAIac8irWnHzl5GoukQ9uSFluQWD/4pXrJ2dIk1k
F+hGahMWeIGDMHFzoZJMVjq15wPdFiWqL0ejRIDXNOlOd+doCUL5ayCoqVJc8JKP
dtOjzY6288ScIKtptcfQS1+SJXP3Gc2svYFjl5g4vyxwba7ZShh0Pqg0STVOgCSU
kFHyu/qwKuP6+vshwcP2JikRwk+QYLqgK45vbX/grFxgmAK33yEgi4tPwGBVjegl
jQDrPSIgz6DR1JA02ajrtqDdJkGuDHBxKFEBNXnd3x7IgtkbH8/OpAztcymeVKC4
6vLGj3E8Nkqz9/7evGTPE+JCYoukC6fxmMqK59PiZHHJ6A33STE3QDFHoJLVBjX9
z5atkcKHEmIS2QCtcxHE+jidUkLvaOeZ9rQyotdBvGmTE/UFre9W8DBY5GnRHHAy
ZZl1jlIbC+lYj8+YoV8HLJig8ZphhnpjvtYR1Icyd5UOvqS1jyT3C+aWG5/8NSAf
dhbrU3MR1cG9GnBMqJ0gw9aavjJsWlp/7UMulx05OuSgJK2G94/VOaG/64eRejGB
UEqE8OfEEO7264aVXFdQdlFLkO5j+rPKEOwzrqIUNsD+pcua+hiMYV6K32gAai3e
WMiHTW50CyYucny309G8WBpY+3DayarCwLnkFKepd/2VJHeBJ38QNq4oCSDupXOs
jhdTgohdX7jpHyGoiQMUurQktYsJyXhVaA6bP33dBK2Tu0hIex8I2LQvJyRnjeEh
R3m01aVUYBRqh7oL0EdJOWcyCGDNWSRmJJYiZkYPa72VtOKJY1qhnys0bL0nnh2R
waR2GMQC844lZlSQ3FfkjHukL1uR79jFnOhQ1Hd2A3/AxO5aohEdxBeCCoTaezsM
6hKeG220ZxTd8U8h/5Ege7xvvsoagVQTPY/CkW7Ng/RQLGe0AUe6/Xdo06MegB1k
Yhuxg7BCs50GeOhU+WkKM+ol74OaxLQzyXCHlTZJsJnv0dTR0jJpFzp31wUdAp4y
xSjARh4dKFIRx7HX3aADuLdykaqfevimI1Hp+1gnxl4W70jLruPsrhnrTg2o12NI
/JPVE++dEp92bpV/aSY/cqKIvro53At8VJPhTsb0LvgzhslyzItw2SQK0cjiMHkb
wNubBz7ka4k97YxDWi9iLa538Z2bKdeBhp0eK1v893FlPdQXJi3DjyEXvWTATM0m
v9AF7uxFALQSAbyR6alYDbxY/fTgQxc1d+lntGiDqGoHVA9D7pLe0VbPf7/mqASN
N4CWybf6H4WfJxgWDuBL/b8hiNLRP4XJjLvwwzWDDfiA2d8QjaGv61dzUSDzPaSz
tLjWIdJHaCoyKH8CsUWFehNCp7iIq+Bazscm/9iojcyYIQXxyot2qv68QUMw4r0+
euNHFjk61Z6VNOuVyLlUIAo+XKzsa9smgvrpEwMovJfleSWbtpyqgmlHTFsMC7z0
StCMvQnzKsRwqnI+6SxJQq/ICjOhUFIL0m5XsInyg6XAAMCDLqb/9Egv0DmHIE3G
F+4Jf9QjMskp9LQnfFl3WY3JV2cWddXJpO5J7b6QVmyDNkAlwWtxKl2z0ezZJfah
2Tc4pZr1C4UmaP0vng+B06/cZihqG/xJJPsjT86kGzzR1VITRXxljwlaXtpt7SIA
eqrN0c0zDcDMh3LIIsvDatEHBcZZ6SCWGi3G0fp3yvgcHJDNX4d0fyAD96YfTtD0
lMSjEa2pLs8R1Lw160HBivGxp7SOOFtirJnVB4EFTlFnWYXi0ujdfbzaFkgrtTyy
BFmNE2w8SpTVtzEfF1YiV6KoerVUsVN/8lBHkFcnUMIa3llU9eJEzAuA0GJnV9Ji
W4FQouyJl4OWQluLSuAIxkrSZKxSCs0J6NUtWOwHsdRFfJvOhKj59UlHNqfPFeen
1dB5XCkf6hNJ7rskx+c96gWj1MrbOy9hp2DxQbYGRmqCqMoDCaJ8MIX/Sv7JH94h
dc8FB7x1yOEVXIv3f/q6kEpFWyvRTisMfOAX4qiuCmxGjSKrSRNoor4EzxrhziWN
TwBvPwGe05AuRS54RnfRVtcPaBzWfQJVN/fd5HqMWMqyTzqaWe71lyENfiNnPZQp
JfUQRODSl+dLPnfsb8dnS6wxEBWKpDPhrOP4MP/JdCFj4L1DA3e/0/O0myFcdsWt
QVt+GwSgLM4DSSOAV4iHu0Fzxtszaaf/CjsddfmOAhIMMO89ek+Q0Y2myLFQJE2i
5cqROruBtBuWEjkiLTdz4SeDUw+W0OxClSuUkpTHvHrxu71DVErED7V7KFEI/9rY
tmQ4hxnEFx2w9WK0xDT862/td+FOl4WIo0ptSi8DrBmHviIJBECZJCRW5A7mJVEu
yRA+M7zxh9qwBHNNi5GUrvrZBfRdlLv3QxBStx8tT+K/24T5QJ66/mfXYNPaylGW
Gmg80gu+1bXTg7e5ztCzgGGUCVNvC9uRdbusSxoSa+3BhPavWCNm1Bougns++ZNk
ZY1V2TAo7rKKBUsUKPtA5lBkQ76jzV/Nw7VQprbJMAgnDTVOoqrhGmVqlpZNWtvx
ryYxs3PpELpGtNPjpA3hkiJDf0mbUWEtuXutR87ImFrB6BSVeBl5csgJV0aXMd6y
ya5HRYx4ywERy9hUXMPmSi0K6QfBFfts6VZTrtR6LS5gPvS2VagNTi12P/56VEIt
DmilbD0OTDfuU6k1Ea56vT62u1aIXq6mBbxoSP6Xu4uQTkciAjccXN6rUIrPFOGS
+aMhQ7iB2797thP5y0jehocL/HEn0WJwf/c4rmvd8Ns5lAoCX5jbYI7/6UKXdPR0
FdCWcyd7TRvZfUq5L0QZWAYSIIIkkRIaD+9qXnEdoBpVeLtgT3hR1Y4CV+yAGEYL
8fX+AWIp9lyydxhgVVmuog2n5fJUfUTIb6kHVwM4lR0N3UDQ6AMJG7s6iz58pRrm
Lype6mxWM4ko7lqW3fzjZS1ugD6GMkL4tIZyDA+SOi9WjlA3egXfQS8NdTSNMsGa
yQFI6aP5G9vPg3Iwq7ixa90NijMwS4kSmxQTuhIVHM29OZgP7HdGq1H0wmRjqge4
LW5XAR+9kfawG8jVs9bYgsq8/9lIWQftUlQYGDMjzXdluIy+85xSjf5Gfbr4cpyI
SDnLshvTz2aCG/aFTaD7OWP2ybvWUxxEQ3ra0AAMcisyUIUwAkXHv9GhtQ+BKxBO
wjnjlgmXixUqaaMoi6IHEFeze1WwrPwxewMntu9FAon0psFKy8M/ykbn4vnx6c0q
Fo1Q/ScVHkLWO9yYRObxTKbCPbmLsjIXi82ofq0JlKKC8EdmXi+nUAO1V7rp6C7T
8gLx9dMnBd7GIT6Zss2BPIngL87ppg9wReNybqwNloNQiKItSv12SKOdcaDXblHs
+rHTy0J1x4qhOlv1Jw7aYqC9prvqnINtiZBq6nqRUJ814bL2KXB8XunkEBLkgwo2
C1LwBfrbS3kFjYKibH3W2NHy5YWN3CVgCWAIyXq/KuEsgzvsv95JnF8PkSYyrvES
PhaV/x2p2/jI42tS0v0G0xXqKVfN29Tl2VBtC2e5nlGVHpKeRTrWnOwadthr2CuE
Dk2dE8y6wInNvpJ8OLP6IipIHe+bOeeVqVNyqgQtSR7kizHXlGsFMX5jig788C57
JGPtek/HxJdZXf8sz37b5+EU+624lZpBQpNMwas5fvy1iW6aG945p5CgaaOuWgIu
J85rPYlaXda4MjUWJ+v4T9da6dpbzCQKZ5YunENpjkAtVfjbXJPab3qZlj7DxWbZ
zCafA/T9snRwrBs3fq6ZzP0sCuOCfCACPG1T5VYBn378v+EepkKmIENHEzE99lKF
9Y5EHFUtYNnyQEqPtZ/GmxsTyWNpVUbv1F00yQm3KYeN04Mmh8cvt6uO/UVFfQ4f
rP8NTwUVmOO2V1Sd8z5RVGerIuQa5L6oxZ/Qa7mLjkFcZiF/OlnyKLn+VPoFMXqp
KRBlKRJR0MDKapJxhllOIuDq/Rzr0zdA2NmE2hqych1b91e7CXODbp9puwNVv4zv
iPT6v2d/q3J0NobJ5GLAh1stuxrp0jfN3JmOgxAqrXFJBVwCLvCRRjfRm1ImkzdS
cilrKdzErPafKXjQG4vXE4nKqvBb8ojnFNu76zMUqmz8DLsrXnSIyKSj2Eao7zKk
Yimcp35EWrEfKUtvgncysUVMHuPz9Xv1ckly8NqYz1VV6k9KpwcY0i7v98V562TO
fB+Wzm5xvn14HC0ZLJuFivFA39EjKq67iLfL+hb37CBBgTUJNOWzliNv1jXjd//r
vA14ItNj5abel4a1tt6GV+2iBGbjr/4yTKCOhiyCJKce3L4EN6hBTzM7lmNgMdcr
foOle7mj+F8ZJJZq0sJxmwFXPWmgihKWD+0G2O4CjRWkFoMn58e9B9YS4Nldz5yp
M6nDYxN7gyGtkGPX1zeH7TbTdSMwC/2SrU/eHzFGq5c1bZAL3h2r3iD14FGMbA33
0XZiDSad9fYdsIKM99NxXbdnIsEgfwMUcOMjwdDNbIRngruU1e1euQfF2TbWynW9
MKi9cDdcmFs2voVw+CZ4zy3y6prEJDqBfuBUz0vwhEYGS8D3x4IzZniKzIbhLDYD
N6BDikFyKD+FSvifRoAslSCnRpYue/DJ8Z8+XRIKjH6l+aFFZAqb8EqNixEIfqfU
V7Uc9tioyJmYLLt+tcrHY/frQ50cj0jTmHWrWLV+S8u4FkgD8vkvCPLmKp6tXqA6
ITJCdExylp9a/wykJllnXXOryHgb31jJI0HcDjIqIJQ9CWWl8o8mASVJ2AkeK4kY
LykhqHhrJFONc5Sd1MR8KOyObaaqqCI3Ku5LsWq9B7nwOU1uplZSwxlQgBa7mkUX
TkrTFMNP53YZjLUsq/dC/wuQyfoZhWsW71dLsXBU2BDJh2/uyl3ZJTXVd7sF1q6t
Mxdi8UPBninA70FovUar3g/yRa9Mf0EH4LGmJNUvs2KmJEIOwEsIYo4Q2zKi3T9X
TaKLEpZN21UtteIyyeDu7W+caoJSHKZqhDWKn0SFLUGDc4z3tUNw18054xNx/mhP
vXHyubT2iPWf2sp9kl3/tqp06WAPT/PVn+EsjJemx/3P99LGQo9x2WhoGMD63x4H
ZISSUqSMNrJwbwXn3XBJlFHCDFifXOl8VrxpMKMD9Cisjccc493FYQ075QFupD8A
R9NNQLRSQ0VTS25xwyWG+bbrdS38Ovvlz7iossDgEdbtSCX+AVgnEwg5s0G45I/g
h70iwacXAISuVJDEyRf/UJSruY9FUds6PJ/4UpTeWxHPI0kU57hjXYLt6bWfEpil
G/ATTDPZW0usvSA0D/jp6P535VUHb8x+6rzQJU9DUOfjA8qCJcnMLXkPINhMJZ7N
N1x+MuLqdS9ezPDUt6VJ1xIfkiAGuHH159PwKS98a81T1YaIhogz2ZYE3U+D3Qgg
mnN+GVMuYPe4I62fccdFmIu/oEIiLabldwsig3nJZg10+4gh8/KSa2cwwqMhGteL
eijTNVZBhFQcsomNAK0A4yFU7J/i4se+bpJK1RH33A8JafaPrXeE+uepJIPIkHjf
GT6Vw3CzMO1MbV5gqPSNMUDZaPzOW7IFc1bixHRXjNnbHfObHZZ8DIIleDyOGRul
DLjHrrggbkv8weCR9MpKwj0XqhpLntxge4hohuyAwVlXbrra+Jl7kmKb4nS0HOWs
WF+FbQHu4LdFQUiUZ76qvbyXowo9m3OZsCrubZy+H7TDlZycz0UcXeOEF+BaamAi
bAr8Z4SIRGyzIPPz9T6+FzK3Hi56WsTYGZAFQgp299NUZSPqrG1JICJpBH09kuFB
8MQWKcq0LHUdRuFMfKDi7A1Szc0d2C3hw3Y7H7votFoatLApGgTxrvuZBdZmNkpp
ElB4hwKS1tKsWiKuzs3JRA==
`pragma protect end_protected
endmodule
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
EhVe+w+MmSbBHmikUgGFixse64AHNyr4ikpP6w+3mTOL9zSykNWn1mwOJyrF/ev6
8Tq+gFdaQSLQXKzR+DbyuyhEKFML8KijPiwudbu6oqmxY7XbEu3nROctevDcLE6O
OHYiXCDVhINg+lHh305C5WmK3NitlNfDRDF9kWPzO2I=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
FiYqESVVIiyD4uUjoEaGmTK0kI03C9iaNdHR3vJdH4VDfDThDt9EBJrvxC5Nw1TC
Lh1wNc3xMnx96B4VURC+gJS5d6TitoR+1rEG5zWfgVCX2vhNT2HpKxoQjLOuTrPy
JvG4yBj4TlWiboUl/7EsLPNO6y3AXB44A8baurCyANg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
X5CY1vlfRU6Nu863DZhFBENeJgwEjnRPkMb2brmDMqwksbPoOndi9/+Q+WOFP+oJ
rdkKmR2bfELw/tAiemaFsoMzNqa4kMuqsnbf8lRZ72bSgjsG8Y/dE/APG5+66Uht
EJgrshWn1ZPXSSOgWx+sN7ckRNZ07oKfbQm7SKq2eOdvlnfsu1O0VOzUA8PCTg8S
5VBgEqnbcfiC4SNijzuvpvyfdANzqX25td4bGevpp8mlxw4wsu1A33CK/Mp7hTzJ
3G1OHWTq2qjHlEmeHuHvYw1z+g6uJPzw34Ua4bq+UMCJvlXM1bYvfB7lSfJ96zdK
byaxat0vR2pDAgTpsnE1QA==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
O4UaQL2ty3jxA/YQ/etWz+6OeepgqNAKY5frXfPpibWFX3oliYYCziB6SKFRMy6g
fJp579B2czrabzJpvc/icQzZ6x46tMzn1ce+zwSkxTzELsx5GekIVxdzRnOwmjh1
lFP2F8kRI5vkHE4h+geU1Hwgqmo88PpkbNrsVIkib9A=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 165696)
`pragma protect data_block
PQven2gUV7WinmAq+I6rh8ClbawIfDKzwIP0QYUO3Ax0glaIZAX1Z/x2PH/UPjXF
QVdCxmc14pcGzkBAqikEugZFh5fzvp67hO7QLJBDZvcQ9cxVcnQcc3DjXD2l1yxl
Ra87E7osMYzuDFfOpjMl1xB4F2zRzo5d0YA3jXZVx6gkp8vg8e5/v4NkasEBTN2x
NGgwJUrwBoerEE4EXGeKvIumDpySlR+v5oOfZciNAKYT7elKmWbqykG6x6VNJTvB
IgdvWlKldQh8aRWOBrdZbqU8uUwe3cYdIIkEI9j0+IFGYfLQNAyqWVfvxACbBpyC
CXahob3bKEJO/84sdiL3hKpsau219ybK2dbDSOXnBM49C4PKUUOHuW2oHb0zFKFv
Czt577uBKwRw4YrrU4PctihGZuuHuCy3WXf7WukpEJDZf6AmyKbXIrpFB52OfcLR
3sWcwiDKi3zI0IYZMNSGeb/W5LACGP96K+9TmH2XebBCjvpFwb4sLABCR/lQlXNy
E5HT3OrUtQmJ0v4fo6JOohzu7FsyLRzLAoy7765Yv0mX9uKFM7XsDxxTeUH6K7EP
S/M4bQ7vBwUf0kXpkkhM2QvQZhRnXn+bc6WKadulUduCOUnf30nW1GyycvLKjvD3
t9ThM74W3xxlftXmToiVTcn4a3Gotx1oCtKeyv/tLda5v6YWC6DHCd8SDw9zbijd
KKmKIzGdI1L4mWedFf+zmrMSzlbTehtjYyyoAb8wHXVg23qFuOrMa03IF6F/cPU6
2Pkaa5hal+7sxOdwFcI2we462T2PH0gB+KImSGCx6Xb4w8n0q/KJv3U+gTuXEli+
iF6MyimjxRL6rP4IoNrPAH1FkN5CYZFHAPwBj3b5nEtQIC8fcbqpN7wUCY0sokuW
UJ0wnoyQgFoQ0HCZ7MK5FAOO9Y0YiXhK39UPc/g00/TqKQhCBij49u1L3K4Sg12U
6IPgKq/iN2UWrgcMeBT9VuPKDi/tS91LNQBylvA3f8m0ghEf/icN4nSQ0sSoAO44
82Qacc1a/FacL3qxzdgsE4bS4YJ+qfmm7V3CdSWcw37ZakD1pSWt9t7nrnF3DuPy
Ixn79Ee3wMH5TIP+s1BtH1TSkgk+3Vn/5IYpgRouj9jrfQXUjw17Am+uJlA5n8Aq
8aMl/n04az2mXpjjy1Y7RdRBD98sAmfrowEqHOxy2wEeq7IpcHyn/9wxS/2rKQai
AvoIuo43sgQEs9u/44dv3NCogJbPA91YJC032L0gJY+4MRuhi6qreY9dZF66k+ys
J/dUfi2Eb9NC6yW/9U9LxS2/1qQHvxU+09d+ucYwwOWFZxDtmI+jWK1qrNBdGRqT
+SKLPwNKcVZTP7yRNyiTSEh13joZTmLwXyKdCvICCoxGNJgAVwAjm/b/wk++e4by
JgY22melL+wo6jpWdoMwBU0jnBuzScR8ZSBPxuy4iDAo0seo02WinvCwa/EYrr4S
G3iwR43POEBC6iSP4YW6i6MOodYNCxG0wlwEcbHTCTkXsCzO8D2Ca8xKPwvBy34p
bwfVDqc1ibAYN6h7B3Cl+Ee0hsqBfwFNqCKRC3y6IO/FsAWmtTHy85JJus8ZMxfV
pliRAK+Kx+NVsrmTK7iYJspeMDWFd4fXSKpgn6tnYHPe91kM3bEka6IdZuLNBS0k
yupJx+okgOjQ9WSdvSUgdntdn3wu2mRXtjPm7qm/dOe2/D/QyX3V/zHJcfOiOo/w
5pM9PoSl3dhEVN8g/AoqKeK7lhP3Xb1zxz91WRBSFEg6JEZvpeuM0d2dWxdvYIpB
AwXKFp27wmP3EUlKjLgbI8J5A68KiMLJHT/IpvweS1QpGU3YjmuNhe5r4oqATIv/
THf2fgyNzo6jmCPWfIcg/pijYBsdeumsYp4hnQjR81MkVCiCGJ+12to8xMop/FZB
I0+Glau3uNe8WfpEtn3yTHfu1p8I2EnT4L71Oov9Cd5icjrhW6cO22UbiOyKyyj/
i+XPPtVf4oLHubiNFUB7dDnWM296ztzcQmthGdKoKa7Qau+MeJNbZE1f3VEvPqyu
XEERZsqxcEu9k8Q2D/3WMkD5MdLoPAfVviGYKesnTHzi0YtOqtq+uTRZDAkKisz2
/OxJK5U3rRYzDRIgMVR2NsfWgBaTslg9uCq38P0lDU8TOFZ4MuPj/z3iAnH1tSOw
kticuZuprC6owGNW/wu3AnOCcHFfJ6pEGpzoziojBAjgIwpTHiXdS0w9t5TNhQXo
h5DkHm49DBogIuFE3h7oNxmLVm7VksDjYnEKTO9WTuOQj46iYUxh5ENpHLArd87d
F/8zXY+TcqFTjNJB7fKgsYeNBsDAL/xe+xcGypkLTCac1D9W6XXIzFLd8A79dwyP
Xmj6ydsm0ChprjrxIKl08VuDxtwzrJPfaFOU+dz9E2tM62MGvP1woD0lJXXXGeHp
xaGeHxNeVoZDrlc9u1ErLr9dgGKCARlZu98aMJJRIoXy0ka7QfFa9HYg/IQ361sY
iaFEhnhUDTEl8HlEdXHT1Gd+fzDvfOT42MHzTyfNeuxCLq0xNINs2z2sFZhTfZ3r
zoqrwlp0S4CC035LM1FqXpkWB2Yu1oOX7J25njvGRVqF+Z5OhVvmdJZl0YGl2/Q0
f41srf2AwEi2YyUB1sLATARWCGDX2Q9EdNKQ13+GBbRR3QCJPdv+ER8TwbyDVrYF
qw82LVu5D2GvvxrC3bdXz+gD46diDpYiI0jR8Id6xE/3dyATD4YpJ8GSzmlTgPUF
Rqax27Ot7xZxaaBHq7D9twiNb4MEHbfSHQP7gxR6Ydj99whx1lu7E2D4Rfc07u4Q
Z0iHWLhC5DFg3rLgyK4YijT/5rMeZgXyAY8glhfD36IpcMBmS8eoF+I/WT1lCpBx
5MjlFH3jHUnisy8ABXIRtgi6NIXYS+hcgt9Ry9vtxmdF1FZO687ucxT5dGXdLYfH
6q9v3zj8CEFwIhBu6U7y3OIW2YcJKk2QwBCyUhJ51aPE0Jy6+AfTfMVEC4zeEkSo
Qa9IcILVnXJj83Qjf4Hveh8Ohd/BhtUxumJMXcUeuZ08kzjpLaOJvnl/v6nS138d
eJtd68jwc6xpQmcoAKX/MqMCYRpY7Z7mDXvUNvM2sefDcM2CrO/QKA/6C2pBRFMm
u+3vGpwbIgY7flrqgD8vYjcQ1HyfT2H/SXOAm7uyZlYm161Eys8cgPWK9O62pEqx
q9ehtCgpAks0jtedlgcqzJytAgpLACDLGGrYX1YW8N/1VyW+OZdE2Cp0rGOSTOzA
jZGGgprkNAq9OJ5QLFlmttCs+VSdU6FfS4QAC9yHqAlczA9pPiONr7aqOhqey4Wg
7H0yHh5mls7Ibi2gGXsdZgXbOUNz5wCmpYwK35bWo+7ujwF9k46n4riSLzFCtP2h
tXsYV8Txb+oMJNBwDCDX+fCc4jWTtct6vwcTYHbpTFK8hhHW5p7xfGN+DYbPqqWu
j1h3Y95AEnyq+yGTNhdlGk4aLUumTT0z3saXQTZdc3gip+p3xW0kplLuZL88r/n9
mjibZ9DOw169MwRx9BHSnZI1Z67KeuNlf8nXZJjnwLZqk5Npgy+hwfPchFWuQzCT
GP8u8udSgTQiu/5jlWBxVR6dEpXcpQN43L39ETbtJjcBatcHBl0ZTN9QRAloEpPf
26YVyw7aDEPZNFYvA38cBd2yva1jDaZoVDwL5HlnJma2UrZq7kEaELBUEuyGR4cq
J8OTfDzwY0em7q7pynpqfGq+0+ifrQ1t3zGuOK2BBU+BYsfQ1WtZ2TtZNKPpVdy6
iKg/lSZ3iY5dnofL/owxTUQL3vqiSD0gUDnZdGMI1kHreCakP6eLAcnJjWJuEB9M
OApMWmyUiM4xt1LtiCKBgRP306gXDUaiSkEs9OHzn15lZEFitXIwB6VenU9Q3+w0
6W+tH5sk1srOFYIcs9/F4edrsQau5Y88tESmnKSIn8Rst/HIlxThISAXQoZpG+Co
+7jPd5Gp9rAcpxEuwmTpPS9rnuvDwhI4gC7gveMQNnKvdgIPrfjiXfxrzY7QBkvR
hZhnEfiRFbO3XaRl0PYbCXEEyuL+rz+hb2cUeKO1PftaWyL+H/S2/u8efrxDuIFy
KcVWIxiPZ/56CjVigCJUtXvQ+N5UP0joBgFmuFcfrQ4yrgl7bClCneocscEuQtet
2+f6mtC6jhra/XKKYGQqwRXVvXxztHYqLS0HWvo7IAWzEeg/fFnMx04NpVy6sxDO
BzZpnyxhppBGMILtvnZuVCG62nIRnJxdkn8fuPsYTVjyAa2e+CZSEojTiHutGl/K
g3DvFNzS5fi4b3cWojSJKOwPZOUlqR7Ztx0b4Ol4RjlGK6wfl14sDruL3RjcSwPO
J/FFmlLzAw7M2HgvfGE+YOu9hEa0vQiPGvn6vDgG7H3waji1cVjGV5NRIdQa6KsO
ORZ1s3rcE437n+Y4G6yxkO9KfXDQleAWrzAqVc2Xas/kJ8P9B9iGyf7OGhU9fqPB
5ac84fyc7KU6xvVR8eNuVZirUuzoE9BmOpY/aEF6ZJjKh3Fd7Y78EV52JvUCO6mi
fS90USRq+O4ivkcVAuNEqWO+n15Ps85Gfq7Pd2MLTyCXB1NuPai5/HbwKfzDLyaY
Rtx164Y5fywK4uoX7m6TSPAb4VlIAijF6MyAMqN+hu/jQ8c36y4oaK4+3Vjiu8XS
E81dUbw9aibbxkrSS5IQqTXN1D9FeBZgXMeC/+eGM5tNWx12EEQhQpbDK5T5Gq5f
g5kjpYZawfR7Bj5vr+VEyffyfa8bPHwTnaDMtWGbIDh+836Ziq5gsmVr6FCQpH5O
tZsgaFqT0TQD/sNPR1hTpMDoXVF0xzQ8yqVSWUFWQhXbjyFoBeeTWHiCmgy7KZfk
VsBy6uxXnH/hjdgvFcYOmFLDozj3fc8bHkePLve7q63LwG2xStdh2bRmjbB3fx4N
oCA9P3/x4ybR5PqsS7hN+AanpOodfHj2TzCMdQSanOXgvNmPDjhwbHHU8hKEkjfV
sYHcUyFG0wrljjH3vc3Kx+5tGO7CHvgoatSRTZw3Htbl85tN4epWg8KjN2PB8A1x
TPRblN26rJBaRIf+BGbdMKfTIXd/rtSSyN/6c9phLi0pBTzxBIGTJfwunFp8BEUx
0DDkYd+0LHLpQBN1RFCMSszYxX6fgEY1OI7rxxAXWqoKdhj6gsmL7ZcwhoEYi1ms
fNauzfhdFORhBbkoJ7TEOagiPpVTf44fMQPYrtoONZzwf2Io3EXa/opS9uWQ8U/s
rKhKbppi2d7IoichYXItfBoR4zEDf5QtpiHWcCTLQTuQgzc3MhQcW/gwPtl4njB6
9roa6smDyZzbl9feKCS+12i3N0mKPmC7msJaAnaDm+wP2o/lMa1yefXzBiPBRSjc
imZYjGvfgsqk5DTOYyncWljS3J3chOvaUb/rBV36CgsfTwEd5zrjFlDtzjhO3dhb
Qur7sOoBChUJdQzvyMBowTPwiXC+zro0oM8bvThqCn8Qw80YK/qYQkz+AF2MsYpi
IyXzj5znnNOzF9dzZ9FMe9AOot7YhFaF6oD6PeKGqP09Os8fr+Af8SktMVX5PLfX
RMJ9HRPuZn3b5WvI3OG+oHiUplYcezHsJ1yL0MnTaLywqD0/k3OToUiEkbBYoTBC
nY3K1ZnhOZFO1owo0GoK6NUH0UtohTaSwtjJO7Ogoq7b2/18SUzW9JPDJVX/pMJo
45yoZANaiHCmfCshFzqDY3dHOc6SvATMDTkOtckXj1Q6KG3QVjWOks8beqGVVWaK
PRs7jvoMJ/S6Mh3vpm78zlRb5Qw89vJwV7YzvCeLrGSjej5ex/9DsR+iENZ/WrNy
0zU1GSD4xIObRQ4Kyg9aLdv4UKAyatyRkVa7b/p7SgE1/6QKI5JgshC1Vxr4nKg/
A3lhgL5nQVEsPRHUOAt2CoyTRhGi1Oc5rKVVLTCPoEPz/iIpDcVkVrUcj3Zmf0Jl
s/Fxte0ntKw6Jx9NiYELFPqY09xksXcdVO+Ls15fpQfFykPEpns17jjA7WpQik2B
b7M/bOdjOlFT/cm9SCf69mhBPTvqarIoypYIUs2liymBLd042ELfqs8uixdmkbo/
LNaqmB31U2J/BFqd71O4Gk49bF11sHlVvvCuGmkPLT/2xLidxXs/7672T40Uq3Lo
fSFWoaru/5iV9/MIpzp0Mvt+iwRAer0lZRUWCuDpM1RqkTzGrOKpb7YIs+E8zcX7
OIRkngS1L5X2E+jIREdcef7At7EgEeRWvoJoYIIhgSFv5J4RW84Ge+IWCRdE7BDt
jpR+HIchwlko3/AWKZy1KOEy1KoN3jZ9XCyKGTIBXI5WYLDlFuAWvNnzQ8WJ+l0P
SyndRzTzp/1/YioOP5dCnQx0QDMhRfpTXgxVMOTqnYtMmrcFfbCfFPk2jrGskiYq
C6+hClqguF7yuJl5AV0phQ9bwuuNOOxfiqBYpebpvmQ2Ff1uzbckSorA+BO5MrUM
92GVRHqJEGs1+AXvhiL+KHmMb9VUZw3tfL2+tj3P/9HJGjAylOc+0aD/Yg263on+
5yyEVuWhzmE5ks9khWC9HgePlKCXBGx+vuFtp1BLencv62Ma0IgXk9t43NnmVSe6
MpAHXdwlF0xD1PLzCD2nkFj6JR+N/saRIhk5ND2VjY3EAQawx7TusCE81uQfUiEL
wnrEMcb0Lzas9Qch2GB/idArX8WMZw4ApVxiAg1xpGNLyPrMfBQOF6376ZNAfSKJ
hp9U7zMFA4J8fzU2EFmuCIQbTpra6cVENmN1ude//SReNOHpXyb5tNUXXFm6YAKb
ffjLJ72+mL/rNNj9Gv+IjGsGos+DrwZ+Y7xEUPYCCshUD8s9PFBrIEKJCC3PsWaN
quupky+S+cAKWB9J9CAoH7U6dDUMgn/ysIsDKORIr2A5Zcxs8I6Dror+qpvSLJW7
ggco/4TH0ZjvhtkjN+mI2WyAngxvQmntZhg9ye54tnMMzqtkj3WAv7uhev61Zo6W
ThNx/hozyaMgapj3RGPKFFCHZLZq5FfM4Gzvq+CmqNs1kD0rHpoBJnOZheMgBvJn
A6l8nnOVrRLQkW5deKZGR+qjIPUoNGfOR1IqYmMfXDYJ4pI3XYUs0C+tp9niL6+J
AxqYkNEb66yp/CYYXhxJYSWp/oYUc35JAL//9uvI+GTytfi1cFE2dcCLsgaspLDN
Qjx4Dvav8EuZDEUWFW5S2jB1j1RgiUWDNnwRWYWwJ/LPuyAsHUDt4FI9kjXYB4ee
Md5ntbGkSrPHeV/xC/AzCqtU90KuxRBKs8iGRuEgeo51rAzmnngs4LqpNEKLp1F0
oSXFqad5Sig/pa66C7O4PlO4aGe+Yh3CeiYDhHSD3aDgJonBU4hs/+2+ETPmROmX
RWPU0gyHV/HGHCCfBaZ9zJ0bmaqXn+VW9CynDS/XMHbBeKWQE04x+fhdKgsimI+v
e0f3V9fm8zDp5DRCMDPZtPvVzcQGkiWWYcxa/OG1JDSxlor3i2a7PWiyiraNUab0
RjZUDK+WSobAz8ziP7+McB+2PZ3tLzIHRdpm6PgCMy0Yy23dsn9QEMQ29YKYk61r
WwVpC5m4dEZaZoo+0jcgaYQ2ujSnjHviB8M25b3tIsBZkkIf8QsLO8IrsLYbfMnY
UWjfxYmHqWCj7ZbStzV7pcm0lfUHeFnikKeO7hFfjMpoZhP0yjQA3HytzNH9nw5R
YY0capPKrg6e6s9oqm2NFSsHbDuXuVb0HK0fRIrJpBB8/72mNWUfeaVEuwfvY7zc
h58F5iAolXMki6Ve8dAGkf+dgAfM1m3IN6dOhXggTkq2H1khhYxmhpHvn9zrNDoU
iNFLF+pdTJo4FIbzfvUMyJux6Y6e4Lx370euEWOAVMycHmZUYBVhiPM0K5f4dlYg
ZlVK7nMlqL6+0jxkA+ItLkTHGLcXF2uZLpxM4GNvj3tyrqdgLFg5Ph3jore2Z8RM
zr39WenSAmbbkSA63ZD2KBjY9sBhzRH07wV/BvaskAt4ggKgkZBQH6Wi2K7ywTGr
BFKUSYi2CMAl8KzEKPDEiizrl/4YZmclAldJCIH5KpI6Abr5WABEqE1wFRpnEEVr
ToISi1NWpFgXqMcGhN6ULPq6i+E5nym4yaHlv+bKRWBRJvPh2vnXv/KQl46dcJ0R
FmGnkolWPTZHuAFoX1OldNJ9MMBVrt4JScZrrlLkQIrzPzwRo5VWyXXhlpEDRZDF
gUAvIumIXqGUptd8QsAfgtB9aLwTAH3M9X0ymaHD/ZkqZJ6jfDO1t1zqnSo89ACV
DW02WoAfoUgo+inpTOcXdJmk1ElUO03TVo12oH2UvZsB8Ww2kxUdGisecWAWwHSS
tB8RXJdOcVsNSRL7Q5+aBOh8m4/d9Fjb0UJ5v2staf1veB5bPUaom80x4vN/WseR
gys8sQaN1IhPnWMARjtJMWMVwFi0U+N/wCyQXEIjDRg+7Kegx2fej9ggsP5M+NRL
5Kj8KuMdzAPhGKQw7AlqA1SB+MzH+s6UTFR8qYww+dZ15BD/c5bLx8QxjDNg6GxL
a/wGN20HK8F/bjACesitm1pM8TUViAR7fwVasrpDD0ciE3GQ6peFNAjpVLjB5RNm
zd3Ul9EgCndvPJQgcuPWYQoYntlFQi/F3qJm1K5582rBYHnY9MPLJF+JxekF7fRi
ujra82xh6UoHc+XiTD0vjWLyF+tyazgVBlMad+IzgIlEEZ+gtrkmBz1TX7+svVlU
oFq8gDljXD5D7xGIPDjIghYMfYGviwSyXfSK6E9zK4hFgcPJ0E+zvNMqX1uZtP4h
qxQDQtXKz/pYN+BdUlAPW6c4KNYW7WTyIXf1OudfPyPv8/XwYaiX2Jzws5Kbmc1Z
KbwqNLBiiwnMG5nK70PwmY7qFLYjNAXd9RKpwL77leMsC6BBACjygAXiwjquy213
Sc1j2iTpw/UFwIyxAYvVU4EkqvyRKu9DrXoyJKe5BhwntpQ9cO7PBpVDPGUBiVpA
lSXlvsU7+HSmISAXomf531OaqKQpAt94OENmK4PHbXf5lbg50O1aeB7KsQLZL8je
JwkgPPtIHYlouud/LGbCW7+ScGSmJtXeCxjNpC/331YL9NeRaGdjV43M7zx94hCx
DLMBXtytsQskg/y1lzUM19MqsoICWNkkK6o123sUZobYMfF6cA2iRXUlO7Z0w9MK
qR8hQEuANsrwSJdK+QaVsSpGEv/v91uvR3BXpvbjdrqbqkWsGGD/pM4+ruey1/mX
gS0Ncjkx8VYMWumnkTyU6n03HSoinAV9JLDZT2f5uLGugnLWyuuJn0mNYMgc/jnY
R0FB6uB81XjaUj5KgqS/INIjEwU3O9A4APVqZEdFxbz2/KLzdngcwzMBbFposa5A
cmtvtTa51p4tNEhfLsgGpZFtmOsGBnE35FRr8OaIbfOSMrHdptSj0BPn/ZHe082x
v870tEDhb/bYH2ZlXumMWOzqvFyHmesO4jGSs8q9FqP8NHlR6v804estybKn/CCg
jHo/nybEhGh0Pnr23cSwkiJQ9QLZOzkFS3Bk72bvEVbFsdWfKJx3c+giCcSBwpQU
Gz6qWo09vbeSfdC4KLMD2eyoiueaP9A3ZKBDHj9GZjPiTmhbT54v50CB7F5QdM/5
ZeFrberPm5OYUsQ0YCVb1S7+m8AGuc3pSUAEtsvd7/yUkLLWMBL2PsAd3e20U/eE
fXKU9IYxBK73klTUFjo77YMoK0n/yvValfAdajymjpJxTvEt+jdx4rHc/osGONOo
9KxXs2FjcomJtM1qfwKRpzxkoWFnPFpWTPOyHTSUoERcZUXFS69mjmSsY3+UDFTT
dFW2TPYlbswG9iTArCAAmmx6h3ZFuzKP04RU3GGbn7m8SKImJkI+G4K0FM1OowOz
ktlfuj3CL06bcf/SHNh8aXb+axfs2IMI8LusZoRKSW8x2aPw3W10B2ft+sa3A6g1
U9y/a+T2YTInFxd6TDNknc2T1mRTzLrvzzHBxl5d7W3vIc9i4hfJxbQO7xrHzBgd
PFMmaZojKz9uNK1EV7AtkXdTJSKqIDLeNtJhL7BWHgnauR9nv+yuoAtTpGDPamZa
oLqxs3Zg+AFiE/Z7iZ9jOwE9o2jLbmGwdxONwNSwWl0Ds/5f42fzXApSz4lvlsgK
gnpYZWWc/rfMa9tSJjJuiZISXot8y/ud4OZsYM0mkxn48nZqm2/UfR5E1syFPxqL
wmFrosUDqD0KFm2OrLnGFIeA+i54Jv+M27qoJdDik62HWGLMT8Sktvir5hWGigJy
n4o1QpmgCRjzyoTdvieVk2zKKH7WFRJ4+lBbo0Cf4qQE97G8uQre382YktSLumhu
n6kT2DzSjaPS6++uJT4Uc3NC3SA4jr76/Dmfa8sUSXcoKuV8Uo4Md5Vg+9EdIerE
4pEn6GyzTytdDPQIcUYTTMZBbKiyKCkBYSufsM4BcrKiYp6/bBb3kHqQFKB7I78s
4LAqz80HBPBWGlt4tUAnKXdxlIfeOi9w881jE2XnCjH44Ro5VXYHhXhC3j0zzP97
nJc7D5USJRQJXrIpXgd1Z2MzOgYEV5DeAxwhFdQSbCWrChVKUcPs4jniPC9RA8Co
WfE+Ao8y1DqLkwjopDIOglhkTqasjoBaIEUNdstsDjE9vQGyV35I4irR6IbFAIuL
/cSvYInYpqx6c9+NLurxJ5GcE/PIPx3fGBk8hnO3yQo3lv5rNE2S3ZKpKXFaxrT8
a39siiMCN5+gaJ9A0VFxGEmOhnYCkmFUf4TKgxIjX5FBzjIKIdyYFoxPiQncdLE8
ZVnKtM6Ydj5lqRHjbkd0Hu49Vbe8Z5CISbbrw45n/gQfPLwnm5xWU6TW7B0Lgl7G
Nwiziz+ji2TPunj+3agGyoq3ZM1uEdHZviebXyP72jipR842ZcAnM+Ev9CmoqzDV
jhF/ssYOC0XXoCocWL8suAnDS1tA1OSSVJVVIAj/B1DIe2mkqfWcgcRoLTKcKufU
jgD5sfd6rhjJKwC/DwaBErt17P+ZAwrbeBwGMk2fVvdj5W5GuF70QTyB9ThcnZVC
gBYjFnlPafvF/6XxDmdp61NAt2dozjxcQz6pPyMEnuaHNLEJ36ukUejTcaPF+skb
sBWdcnFz3rV2y/qKZAD2OJGeOtxNhBtqBRmW5txTyoJnD0pEJXi7p7unGS131WL7
ANnFADdiqApxgLv+BNKo0gsOaLBKaaRFt8bHvB/olN6ZNVlkP4MykC/Z6BWD4yp8
i96VQ27FmuI7zdE2GGj6GXPnP73QbSUFE4ZA2Gt1uhMvR7jsf2qx6CtoMq7BqtEf
s5chnCFtUM9TSejn5Hu81qMd8OhHgt/pkRQ55QtyVj48oLpri4No3e59j8KCuqOC
pAO8vgz4E49fQPmAei+DFatcodDl6r6A8hj1dcfc0+KNECCBvLbq3XgQuOL1wqTM
d7l/ze/N4lZGhmNsncWamRSiCStNPidcniYpvFdYWs5NxyoU0JJmqUsCS/cWi6te
vcqcnDGi0YStG/iWfVN6uNiS2JmGy8VBMBo2q5jn07wT/+RRycf3geoZcM6pkY5G
JSvaKRpNhltSsA8tYPptkHnTYCibRSun7tarPnwLCvtIsz+pK0PeysrzW+YmP7oF
hhbzXvJCGrwZrqpvVUw1R4l1ZsyZ7i83IBwow37hnS1GaPMlTIMVhZCbkzTVv5r8
OgkjF0L6MBkk8okZsyLMFbsyR8endgecmP8fil9jopYD/XpyY1bgwOxyjygRh8QO
1vkDTiT8T2d1rvBbs0RmIuRomfI6xAOPgnckPFwJyOwwRFhiNq4SV2VxNuXE3daJ
3hUY4cCTG1KvdLryoOapJ08LAZkm9WPSjiudn72s5ibUs/cCbLOL4qB108pciBRC
padQr3+SruJn+0GEvk5nt6FYAYBL65Stk8nRwC0Bm2tTxggr4OuLjNYDhkpbIECk
IsyNa67W6NW+oayP2uk4DI1vEwyaoJaPC1L0Sh4aglXh8Al9Lhp4sgW2mNwln6Tl
YfU0skbeqLerhPn2XhN62yMTRSn1UPUpBL/9wTde1ZnL9GL+o/vp0GyYJ8GJ3J6H
3SaANtEJhs0JYPDE8tS6KYYMvUdGJI84Wfpp34Ah2AlQJlUvL83Xi3tP45i6uN/H
D3nKWoAO4s5TDHp+QHiKDF7lhTOKWMaQmo/h8fe613u9K1AGRKvPbIWUyH2gZVSf
af4x5m1ZxQhPUu9hP8Rv0USNO9+hGSjIBJTguMtfk699HdBgtGJqzIZccOBnKS8d
3+SQ0XG4VKYsiQ+7NkJL6uDpzMmbfxBMl+JirUH/zhKqeVwOZXU9Jq8rM4tGjoc6
4uVXaDwD7aCTsc+/7ZchDRg1uLQhwZKsB5ntX74we1UNzL2/EytedFjkE2WnpeOg
1aX9exdxwcInc/ubmgZvZlm3uJ8oePCdMP8jlCmubsx3dWleU2gO36Q4y9q4kcEK
xO3dAB0qKi42ADafsbLrp/oy3odlICBahl86Bgg9+DGReQZiDYNOzUs9ubACvdtc
H1L/vnZfp4H+SZH8OOPuY1M+3ICOcN1e+pOg8jL1Nr8Cxyd/f9h6tJmUmwdN6DAZ
oqW5KrNhVJj1W70kdFugqPHJgvf2jOLbYRg1lSZNP+ElrNd93xsh8aXsmycDVu/s
gEMtZrtTdrEUo5D5T5PcIa3uQt082NJ4SDSvecTzSLOl4MrRvFxKi/8XjjVElElQ
yELGMN4mRTeTfEn/GKKFJcu60Vuw7JkD6OcNyTJCs3zomkAAT4keYv4yyxXqP5Gk
WxNJm+JtrZgUSdfrWzJGP6FNjAmM/tgJUsxsx64efEnln6gE1PCH55cOwSKBkNLM
di6mIisnxCiwQgOsKbTQLIHtqpucRcYULY1RSiaTdbaixy98lX4io/uwzmbFXWKl
AYt9jgimbEXwDDl/lFzqMeoYGozDyiGVowD/68ZC3bhWLn/LVkNDY4y8wqphgBCg
GIK/pZ4xbAt3rX+j1BnEPLcU+s9ziMlv1MglmcIQ7qntCFpmAQR+iU4Su3WqkTX3
jw0JTKmrwHKGJdWFgMte/ev91E1kDIf5K4pbLEwaRcsLE3zoYEDEM+jQUzxIXrZP
/ydbMKqDowCQnwbw+sy52wACNkm6hl+L9E5scPghhmqrZsaOyMJYyZdFR8f0s5q3
V4TvL0+93dzPoInSvsQfNeJUpVB+0KbvD4Z38ZAG4yCBSCDovL+RVuflI85XqhJt
JI8EwnglFAbxvxe1prXqKrxyYWZXwLainMn1fR/R735dIGJu0zVbG9705eK1SQ4i
d3aZn7DhKvyFe++1J8so5AkSnuuhPGvvlnXXJR4BckzXEUa5HkPgkOm6kpgBM1g9
q6qQNu7PClngnoz/JrdNSnnMl2yDvpk2T+TYtQM4hirfWhlx9vNdaRjic/xsVxZo
zJH0N4JgvDEB590QVUDI0ZgiT1/iQAm5EPa6tTVdUQA9HQUHQHzUiFGKd78aKDV4
kiyxglPRzKNmcdLtvKqtf5voFKdbQC7YaERG3XQHvDWRBZHsrvc6nIkR/+Gcj4Z+
ktOL30WqlAZaYuaMjuDDSTylNSo8pp8hspr9ziNjPNc41Lj51m8s5b/HCbvn3GG7
AxUOpLJeWEeMLrCeKLAfAsIBc7tEFOCedCpr/tpJQCqQF1ekwGFnulnw3HxQOTGF
N9tXUXArRbTcuxio4lso3FGJ32j1zyAyov9v4HCphWB8gJNlkYEoijWnZWrOJJbc
ERgNNpAYRN1rnaUuNhi8eDJ3MLy4FWSch3JOChaM9itcXPH3YU5r5bLuufyneIlE
CJoDsHk8SrviZJswbhHjADmCz5qKUOi83kBfbAs1+R/nLUhlfHHZiSMPhY2eTn3/
JX2/w0A2AsPueL+/q6CdWFEm8mx6FFBaWtUwNt8VbPEkqLmN839QN5TkR1U1edTX
USUgXbUq1y5ToIkPserO5+gE7QHOMWoKVW1e04OnlSee2WsubQ40OX4SaWa3Cpz3
2LoD25MQxM5Ugd5eK+hWs65tCFZxl8wVCyzzYXkmGKoQLcNNjXmGV2LWucqSmbUz
99F9J/8QInvsLgLkUqvv9p/H4HZ9crA4k97Kn63aA5WGTIebUkVyZMu5k6x+Mul5
e9KG8S3kAMcE4iJzGym3YRZs6UDzeVFM8V4y0qbGIhiioR020TJ/fLq6OZ1NSNtf
OggPs55ihqgFdPutOGBq0EWrogqG5OiN6oeFxQKG/Z0/smXOuroQfLlYDiD0/V6v
LkjoFHOCgC+RslI47ImJQCkXVU+54y2HmlE+Q79U7ET1jay8+UMl+tC52vtB8sbU
7iXx40hcxoRL2ROlGAf3V/3aNxjqCnj2hmIP3Mi/JUFThY5b94Jup01Rft6oP3KO
q/J4tdCgIEAnVvTmcA/MBgJRqQas35GQd5W10WrnWb5rIVg68H7W9kg5saHons/y
n6nKtBQwqz8BtuX1efy5+/hY9C7tApffBFMub032AnkZPCufXYTlJcr0uO+nBSmy
Ie4m5csCY1DwaP/wDi8KjGmHYCJcilRNEz8vK0/m5KjbaO8YiovmfEbN+v3c5jVM
ZwLTt+5yWEWoTNwI92bR1dOngRMeJf8JIGmUmB+n1XN82SAgiug7tXOY2HjEVu+H
HR3B83vxbwwdhr3q8lJLzo1cgCoj5jdwz3Wau9B9hEmwFYvizDTshI21i8YqWU4u
7BRNu1dc6WgoXU6u0WG3RICb1JCugYezfn9Sbx1ZTBZyw6o0nQbAmnkT77mdOB44
DgOH3Bu76cAtfxILOGfa+8JKn6FWT3uIOiDvdvQV5bvb4EhyCaHGM3OC4sOy2XbX
0ylNix1Rla1AdeAq+Z7Pjk0xi1E7MjDYUGNqYPCrIqTUUwgWRmAPtvBWMPi9AyXt
GyV90GpM9xIWS/KH/mPSUIoYEIF3urrIKeh9Aa6Ew6g97iVmfFoPd8V+cllA+o70
hOKONmZ7BVmX+T8bv8NsUWRXOtK3XQzJbBt+1r+AxdjiISFo2j/0VOqdwmX0ywiT
jj503IkOH7YBRuhgB72nICQjBxYDBwZckg3oXrRDhzhIYtUjua5FnPyITPh9+BFQ
xJR33rQ8Z+XjaJD1CkcUNnnA1qMmEbVZrd1MY1gUaGsGNXHgWq09AccVjU4XjUJP
0hcjMdx4ZzOaww3lDqij2nIZ2qHT0EavHu8gh5T20E/4vHWKtDNyG6eUsXjcUvqE
fERmUv91wYDImvKOs2TJQcYYORUUWGiCQO1jPptvD/+RogNMncA/PLEATmotJXZu
4U5uS3w2C736SvyvKdRW67g6lucewgzQDShyYYN0hqWMVMGi/Hkyq+XbOFgHJZpI
f2u9L+8EhJ3V0wJunIUeWPH897PaQ+8E+6mnT+9m1FgQ5Sf4+fugU7aNYDYJXujh
uvnTv0m7YH2CZ0/MHTR7yhKQ58UGhvHQJ6ayB4oLeHMFjniLtFGy83/vWVHHMXC1
sehBSSavBfhEWs99QUfwMBrLp9EdP7aYqoZK0bRCFWlrba7l2LQQxCVd6Wpu8LSc
Hxn1TiHRe1CvxZQ1kRBLIZQ7A5ldEH8qNtrjQYu+zSoZE/TLnzCKW5RRjGuqymQe
ppqR9Hwkx1gkKfYfkIOmrjZFVmhZtoaYAhVgbtD2yDAvC+xgCguhfOveonuZqqMh
BQPG9sf5n6IEAebbwZMTYEgFAbtjJ4RSX8v6X04i+cp3FsFPWX7B5GjZv1BrBWMI
C9ziKV9rGASS3Aitejh7TM1zOe7/dgLpXwgCCUOSC+vPENo0on+fQix60L9I/P2J
Rimp1Eq8Gg5tcQ6NbluFb5Ae/vWdWKfXv3J8z19MmdhNP+Bf+2hMvheLhsQtrzi2
Bv6c43JLUR4v4v709Af9Hw+EmNHEVXYkIpguCJCEElFVlnVATf78F62MQ01GAyD9
VCo/FAWpOXaEPaHSqzD8Hmbm1xeJLAqCkQ0YqiBPQoVKpia9L5h0H9hTP8kGl2GY
aHE1hyq5N0oI7SLSV/lLLN3DBlc3hqVFAOnKhmA2zm6llBZuv1N++pqGAOW85mPm
TbXW+9eZtUP8lZZJ0lhptR69X0stlwQe8r8MDcaq6cD0QE17O87Oa9pa2t37+0t2
lHKV/1KSuxo+JH/K8xNaWwu4PzlEfY2PU8soaHn5CK4nSU6Ta8E6pzt9i/lIIJX+
xoKRnf9ozwYPvsB22KswT6ZrjmChbfIH9rZRIuLKmQjHZCLvuL4Ek1Jex+S2Z/HE
goMGSEpeCRZ4eQAT0IZ2zLmEqR46yyPp0OqT2gACAvrL41y0ehCdaK8FDrxse83Y
/u1MlXJdseU91cTLHAPE9GChKX/15mQhf+vkN+5PfYMEUEYkhZKAsVpakbDLQJll
FMeT/ToX9qKJ+hO+E0FNTtKae54f8+Uao6EK3yDPuab3ZFzk5WZDCPlHBkja+upr
0pNgUKNWG49pHWkPOW/YnJsBakWVTDo2TyNE9ooYbfDjTcQrDFgQVR4kofy2xXkS
LcSLJsxKlEqNDtJy9YTVOQUAuKGESQ1qQ48IxQqFOTmDLVhU4a1ODaziNzA2q016
cr6sxxUCLBTOGlTJI6qR4PmwuJrn4kgB55Bmd/H1TbUTAFmib0U6nPOai5qjqxbM
zgT3vneRk5evrEngXftGBoGbqlLw7vrqlhM+dfz3UvTqAvfih8x8FhjNDLkyPK6p
oUcFPduOzbvjZjUUGhJxOJAM6ZjLsO9B0Jdny7QXVvaexp6dk2ZhKFRzJiS5S9ZN
xqZjQqxiZHHX+ZaCdj8HWKL1cfSuhvqw4rWov5uoYhifqpZwlO6QHTQ3n7bMAYgg
/+e6sReFnArUsG2GEav+cxcPl4XEqdYsUVzMYO2rJ6IpCILDLORJulJPg2FqZD8l
ywJxtop04jbtad8H8CWfVY5cgd1HbCAh0cpnuGEtPvn3KnEOIIL2x+NcFOFjBCNi
fTQkApzB5UBIZe+S+mXHS4ZFphNAcZBtKWPBzVo2g/ADzZdu7eADU6ZGMSnPxtxJ
Jp7yXoYQIxjAC4LtLOUS+mG1/ccPG4NHwz+ZYPaenJ8WEQk8OLCqFD0CM0+VGlDQ
YuHyEkpYrxQJasXuDtfnXIrTisuKEkzQAvhwFLsktmM9tnO1bN3Uce0dlR9//eWZ
LkHUgd/BUftOTC3OE9rnaKcjlPLiWuDp4JOCkMfx/ExW1n9HZ4FskQwuJYVeGKEg
1y2gntO9grLixp/cxfw3rXbRZ7YmXcoJI6xUChaju4RHZbVMhxTzBj8yOfFdeAUY
xX11Rg0s0Gs8ay3x7H2a8Uqg4RqMZH6APJd9MWCvjl7Gz8p4EtmAyJ+Y++F4HvTI
DFXFURn0BxD+OzA7fmpHZ2WjjsZftPuTFlnX0X9aa6tPs1TM5bTVkGxILZGMhQZf
JVnlpNn9sAWh+TwQ3Y43xsCq3wA6Ed/7sRxtYMEYQOCQb4XbVv55B6IkGgFEZtaA
bajDgRVW2ubtGYAs5R0qwCnyAdFf3+Gxm71HG09Xx0sgA8MULCobEm3FM+hSUjCT
13KJL5Em7QVQCXzcd05yj4Ka2yz4tgSM7vJ6vmHOqPq3xW+ZZh1tUkXDG1/XjYzy
rN81Z74JUlslnZaBTHhj9KSU6YbiE/Go6UW4qWQBfF7xSXzEDHU3X4APXw9//+uJ
92bu41gNyKAExwzDLIvo1uqdmVI4HbNCwAZ61opygVAb0vy6cVkKrFyk27cgJ4wR
Md0f2ySvByXt4ewx66GCk2LvLseBW/ChOkhIf7bCKqYCfpfd5k6J/WNbjguXEI5B
LFedUjeb8+E0DQXUvwoT2jMkfP5D9JTANaLnFkBsvyVHgKO5jklPDJSH8IhJ9RSe
HPQ5Jsi6uMKTxPlAwqnbc5MoVW2ku7FKPimGCDYBkq8a/V+G354AIAuNQUTsPrF8
WsIglCduhbkuW1HFqKKQE34X4n8LIfdjgyUsSD6qS0VHKyWscBgKe7A/doBGlXco
MkCGnBF95JKEfc4+Uo58PTilmUURzm/B9TZCZKIinivTAacAiZZUCPcQVhR1r5SW
he8fcPOKhQGVe0qbWa6lOeRA55xGOlaWNz9Hf3OvmKLJ/aPhy8/X+Aw4nU/Q+9CU
jqPMHKVbmakAuik1QW1xJtzTMzJ+L6/U7nZVOfSdR2Sx8cC9Z1+J2R0XcecUbbCV
zTSs7IJiXTkZX27TP9V+47iGrt3usFRUDG5oNVW47BWZrb2ZL6z92MCrVoxfUIeN
QU9oaZ63vXTVgOXLrhS/bbhOyuKtJ/IcjQLTET9k4D0RfoJeIUvdEuZhnv8Yk8Mj
UHXjLOFTePhFukHUnS8SzI+/Rk7W+I7BKJK9DnTpzDcZV5OBMvIerCmHEBf19FsC
VVstqIFjKhxE3CJa+0BPcuNXFkXvo6MRF19LpntfkKCAirmRY3hjA3FZ/CF6BG3t
MEhK5oBm3aCgGj38wQtsHAtBAiKn4mGHxsQhq51LN8V8fnkL58RdIj8wND5wzZj6
oYSUiUrdC1QsKEEu2jCNMkT3/8FXzyYgnwy4DzWQDTCkFW0HWtKjNZ/bcAZiV/eH
DOEt+nNn4ARvv3tI8RukRfpx6BOw/vMGTMCOGhUHqeoKeXTsluYC9G7ntFU06yHv
wbw9mpOERQB+4lgtj0H8IY519QG4oUyd69HtjAyIDrk4m7rGXHvYfUCy17CI0Xlp
/RgI32t1YYiFlpPmbCSLeFysVqqc8L4u/Hk5tQWjmcW1N05fY7LvXjBkpf6ZxY4Q
I/nvf8d1WnRTdyunD+GUDwj8Ys1EJIHY16XW5sCu2kR6arTwcaGNMJemThanfDNl
jQ5kqqA6qnHGAptxGDWUmWdvnDBCMfJvpu1bYkHEOM/l7dgmtcsIFxOxCQ+IrgD7
1WWpIxAm40tELmcvywyFsVfUKdHx8Uxhpz2lTpk00g8YgXd/BfiNV7kjsAyutG2+
BumZem9ZODbvaIHmKCSce270JsR871qqcVg7tmE05rKw3dfxM1rZBmlnSzLP08CW
F1xQ8n3BO3ToO8lOQhYMzMS5otbXZgqpjjhpSz4lcVrz1J8fmcB0gE+K6Nbs92pr
9D24utLoAEy2JkldDwcIKNfbbdcsSnacb7y0sb8GdnkkGva+7cXf+0F7kO5JoHbi
40SlwGQvUorABC1dF8G4KNc2b/rC7ZA3WVaR1GNYKQ2gZfehg0yh0cfFBHxiBx8a
KyDrx7pQ7KCrvwa6PIcdESfM19uNapJTSDyx/utMy5huh7BgJlwJ9YBEHsIA1PjH
WzawLw9Cf+bU+ODH2fWDdKYR7x0hbC1JXyInriVDRbaC7Q9hrZCSEriyebWDlc5f
yI4fTDOJm51XHbMxmbtYDoZ18vFYNds8VUeiS0V7Lp3e07H+nVReew+RhVBYXI9r
OqHSn1D9RrjEqMTzfIGSplgzdagKdlP4il2j/C1Nfkf9aPHTxmCMUfJILfLmAE/M
G1/TcBJXJamIz6xvYwDO/5eBxUkttVaNUjX5f2EJQTJiEqAfMgKi4Ys5GBF7/TIZ
J/n8p6HZYL3o6tGM07cTNnZbpPs+E/znmZcTTvSuuPx09+8gXKhuPuZz6ql0yrO2
qTdkuWsFNbcQPRiROu4i0kWKxAmPM4OieqKHvnfRzBOlQLxarlNRVMjgrYi8h69u
MqtaLFQHTx4sQaD6QJ6l9ZXsHVxU9nHRxXgdb399dirlVDPzdD3bHvMtdUaMMjv+
DYchq1u6S5DwqrKUTlPDRAwbM5X4fdC9H0v/EnErWdN0A/KKMD8YydDRZvMwvW95
x81/WuF9qkkXiYN9fSLpcIeAALN8fCdlxH5MlaAAqTnYGtowUxvBEmLRwUn35FeO
4WM7cQMkJXzPe79PJwwsOcHK4VsjTOqvdIjnRF3Y46v2I91vdkdO7lcOTJcE2u/G
/D8lWb1AjZT2k8StVEPhqmZC1kzPtEdP5ZuCi/DxbnGiZ4VyKFANDkj7uNLBH/rh
zHvzvhxTXZq4lkn/WtQhuPeyrbD5Ybwy7v83T3eJd1VTpa20YUwKNdPlvbJqN2ex
W2YnBNGUHJpf//CIWAJaTk9rAuBlGlB/a5oBqdig7TVeaWo6+a58UUXAMOUiFp3Y
HKR7njspAmg2d3Wj+tFvStB6H3VXO+zXdYGuILemnkdE4jrgaI3MSEqVXGO2Gi5/
HUgPGQAucJle+4LmMWR6XzVseA+o8qi+tDt8YdV6Ephq6ibgnF8gX8dmixo++CiF
VwMnFV5sYC+6gXfryEMt2DDZQnx7kzOlPkhCOndCmrddpFSIfReZHFkjK7Fh1vk7
m+sVUdTacRmhClc53KDtTIDgCFonARI0ZxDXYm5170lDU+4QwmFMjF1ItU9NgH+3
bih5lS9i3AuPWhoBjUTlR/Xx+XETX4jtmPFJZxvbAwN2iCaWtKOyeeP3TtRsW7Mm
SV/YG9uOr4wzk6RjjC3pCbCzK0qt0I3SvoHHA/jxjKZzqJLuIboWn1bZkSM/PZKX
5cju27ALZQzC7fPrtSqZJGZvHJySPAdSWMSy/wdu41feB9yRPJcscSeo7uI8YpRx
aCRFI6lX+ljfQpBoK4Hm22/kSAg7XuZUI4lGVU3bZthEqPuZAs+Y4UeyNz+BGbka
LH1Yif5UQ6u478Q/Xfpj/Dyz/eUB38ZVIOX8fdg1zck65w8EB45C+t2iQfX4qWdM
GVvNPgd6FgVr+yxCPzQJUuxbX7ps5mL/ItPwkKpR3DbwZf57QK2YMl7s2ZAmrFPB
9c7fm7DeKa7cbSthnjGg265YF9oy/mfuhLSwIThnkbsevXAdZGVlMhyTXjykEFkf
GYW0Cao4PwkSklepJak3sny6285H9Msf2eG3AV61JCTYn/2V9Kqw6nbSkt200l2F
Z4lUTqbJDlPTtjBVw7ZzM0L/3Gz9M7bu8Qf+sqPTu+yq5nyD95Kl+INU62XcG9/d
zRFVtpCGxNzdCUjBtTkNMr49RYqETXb2zp0ZiKnzcyK1ParcgFu+KOiOxF9EjHyh
UmM17t0qIj/H3ysqQejbruhxlRWqhMQd8y1SaA9JqLdGPBDHJCp0jWokgeRpwQ1l
7cDJO5YRweGoorwv+2LGhpwxtMAGLGu8xfiK78wLvdAO/DL7BcGpHpc6ed5a0fPf
Xkti8pkSw1qg1auhwGTnfxL4fIn7iRpPJEY9exPegyfK+vnuYLQqF403EpJ+GQxw
rZ1w3LaBjGnvMzW0Dmnn4ZB9IyLoIk+zD/QECWEmIVma7bfXmxDXMhp9WRlq1sk1
aC0yIV81ZwsD21ZnPpEGFt3tUZiYflMwD8rty9ZzvrzcdDwmw/6qf22qMGJrUx7V
e1t5FJnn28EGcNkTk8NQHXRrN4tSxkLi63WVTXrXagEpVQMShtuFkO0IfAxforUM
goiQAAjbTqXmEbr+lzZz5u/8SVQxWn2Ti4mPZazEaOQmbrLBz4Lv23AkVB+SFowY
PjhbgyVxMNnASTAxgpluzDhMQvqUWSqoA68tdt314iqpPp8tTlPYLRIDCJxj3/rK
v3qIHW5OrfJxSFjsBHB0jEI/gvV71NDY+N4+3GPFPYSHUVOYTT844SVEmy3Klw3f
irJwZT7geFG4xkSbZQ/57pNH8+BGxG3O42GfvZGFUFOW/tzA1obzYcTuLZa7dSsc
NnbGDFQKKm5wl36q7zzrUOvjD+jKo8FaXXZOlxBXRFLmxFvTNnmhJXdRTIpM5kXZ
MhJbi+BqdXDeJfmJjknEpG3PdXZPWH4Z+xVM3hKN+xixz9CLQnygwWGn85vkoSSw
M1Cj1VnoBvFhRQixxqY3rwoFxKmBMmwkXitba639kKXEUiHXuaQapm2E9+8DMUDD
QM/44n6CV43YNOxxzErOhyNowonW9+Y+dzX40DkTAuZCL14aJByjeR9Cfg3ioEIT
5d7LEmVVale/dmA9f8a11Wh5sacaSKiCuZC10bwqAJQOpVk2GfE/UpfwVeNEGBWN
esJO04A10hF1KZcpkz4Zcyb3HNvM5c1+fyVYhvmdtSj662BdHRwQR0ufADMZ2y7r
MQSiVkEpMCjNv4oZ833NFi+h9U4bBRMtq587DSjS9xB9G9tys8JT4sEYQmJrxrj7
hSTLRUA1XBLb/DP88dGMOoFOumGYFuJolgT/vBYa+bTVCRv6+Gr0BAHTaCuLhPrI
GU3IC8t4gwBfg84G+cuwARX3iTYUQWMh0qFBTcaLdVrY7PykKW4adcCquKmha9Hh
unH5Y32f+JuZlXXuF2J/4q2+Gzc74aeHvZNagd0IvuyWoupHfjs2JJ5a2EJviblQ
QDwPA4fEu3OcqjxTRZMQXJZSX98HC/qk5eBhIzaqXBx8j9mdlNEN0UcHW/9lpbxZ
dUPQisCiwau+5CuzPDUgqtM2nQLprTzwMmDQtLta8DwVkPRuVXvgdJl+ItAWiG1P
Cl3QbidPgk0nHZyr/+yh4iSeDjDhb5qhkNfK3yeRb6QXsgJ7687FuJW6N2AolSRq
2gwURlbhjhwxbBiF5s1OoFIBfrohFLpGUQ1tx03xY7L1I0noc0gQRB2R5VA8uOEP
LoYpwMzJooxRWRfeC7QdDbxbMHQaHm3Y1qe+UbfdF3yGG96r+XNpoo4ayUlCxpk/
hEIg4oyBAWJ5iK9TXRDyiu1h4saHrEJp8bBqkPwDhP76bfZRlGvBFD3H96rbY7Dx
1Mc7S2SimM6Y4GOuqBwO1HtEIfo9ZFMxIujhDJi/JI2VHSjmmy9Wz6ce9RQ4N1kf
rwgB4A1AWDdqsrpvLlX+6O8xfDe+o8je96VzIyp5yQzW7Vo5Eva4eHztfOtxyp8U
mVP+waNIqNWXTnOElpOXP6aySFGA4mdXEm6ajsd1YRSrOYP/bpLxhIpsE8h8kw9J
2uFox3CJqrqh3BTEWi7WiqAFv29y6IKrgyWt2yFgDE1Y5wB4jysmmA44KeP/gtjL
9zWoeqkp/bB0jmVsXp2jVEImEq1x7kfIESt9DJj+W5MeDHZes5nquwHlTt1FV6Yx
8lbHi+kUNU04DZXBPVG2vpxj3fwqj4U8usR9+iCBQA+/yUe/MesMWR11hiCZNS+x
1KFgnYhtjXoHVBmGm7ZYmte7Zeyl7hf9DOmqP5VQzU+7CPltgFXPmekMhL4fQD92
rUPoOuqhwn/NgfsmAn2re+BwQnHrsxEGD9ylJ0z8sdEjSypYsRl4ltyHFD/0bvY3
tNPbJSDZjHNI5reCk9GHKZ18U/AGSdiac0gk5idbrZuXafoKc0G7mNy0CWPHxooo
s+xpwvwaadI1p22JumSY1Su+WMYjMnvRUEaOK/p13o2g/qk/HaOF6CHNy3nMackV
uLy5bJW8l8X5BOB4147lCOmc9nyD+pe0plRGMxqSEiZVK6dlfSY5A0s93tZn5hQP
K9KOxLhivx+fqyM/4/6ixPKoLGyjVMZ0P23bv7mGRA3LgGvFippaOK8RdXdOI5kh
0wzuXeRYIZ1cFjBHt/SGgqDWbVrLO9+CiaifPPfWYT/8dWmxY/dOP2fuZBYHkQYt
wBt+XdVR/90tuc8y+PXLJY8GCjADn9C5zD6m0EFiGD6/Jt1D/JumN+GhM/QUlQUj
aFVq6Z3IQMMqurEw4xbL6XsruEHAtj4H2e207mP4BY4DrzEVZ4+wI143N4iT1h3x
gzKv5c5XsY0FZcT0pbOhrXWviji34Hvr1lLXUQr0PcLS69qWfLRr4DRAjLnEbQha
48qgLvmcb08cU2h+IsCq1ZX0IVtQwRtMP0JnaI21ahVnkAHKV8KYRIVRa7AaQ36e
b1ts3xFgjsUPHLcmbj7f6WaNeutLfJl6Jpjcnm/t07vKyQd5zjmGbb7mWr66ZSib
fVy7mz6ee0NgvWVuNJb/WzEbOJlAwrykLYy6uwp9Kwj6wVkMt2Q0L+EDbOj0R0wN
W7z9TqbAZtHAipgYeT/6rHe+ipQyl7fH2R3fqwp3LPyxYHEGJeDxYfDFckovJNwx
3qkqXGb6LDVtzb1jhWpIF4iM9kcGf/7WVJo5hGndbN1d3uWFIt/3qjaewSC0r8dC
Ur/d1n3liyS1/f4MSvjyqnoag6qE71jUTXvtj1EoSBF+AwuP4mOz+9dP9xnaNwLm
/aN11Dkho8u27UFHl+PNeKhhViJ8Qh/qPLsV2EA4NVrOh6qDDt1kDVkgzS6A/FzR
9A+PzWyvBbVg65bowPWG4dQdgRxuyVn4zGzq3xTO6amuv4AeR4a/vQb/lzRCHzAH
IR1ZvkqAJLqa4iHLabUKdzNS9aPhNjQYlMDvsig00WKURePTseW84SGfReQ24AXF
xNZUmlFDg6uFCOQsi76kaACSOCDRfk7gl6MtLsH0KT+1UQ+qRhf0v9nscgjA/yEo
cl4sBlhw2cfZIYlvfKug1kMqK9xAtGqkEBqnEFEUoocsaOCbyR/tn4VE+66+6Rhr
NKA/ujJ6jb7JKh4PyYkZqS3PkJmz7b3sLbIY2SBL60nxMIA769qjpWLC3NFogAm3
B2F3CVrnOJ0Hri1ly0qEcHXYQvb8nCgYJB+GfIFDVqZkdUJYotTEs2jNX6lazVC0
0/d1yZYM7pOHLjLzOKEsY7J0OSghlfJVCWzomMs5Bt1KuIl/hzfK49uT0/5I7hn/
6PIkYIu4dGc5HHc8pIPEmUNgNuMyQIpCqqCShfMosR8wXQGPPgmT33B3YLgUHNZ2
Ck8QsdgEMH3VhW/8o8ZOxG3a1P6BW4vlsACX0iDK4xu+Tpgpk4CvNpU1+NzrH4zm
VWDgSMHgLzfzq+lSvaEB+Ik3g+35tTTfbOvdMFj4cTHtXhXqmrhevJ8ophmFxyTJ
erpYz9wYo7W76GC3mNQxMZtGB3AoMcUwOp0KRmyC7SJvkFGaP1W6S4AyrZtlPerx
RNTiAXLSbIv/W7KP3rNVEL0cJCj9WnuttYHJ5EL3Qngf42nmfGcLz+W37R6NHhyZ
GNfuwl96RpdjIiA7SR2brwUPJHHsVmwg4qXaIBJad/tqdZc5prPkJ1Ya1zc5NktA
Am5GHK12PBLZCtCcgQvM0mXuMyFg48efttaQD0k4zjVqTxpSUwnGGj3leoqyZek4
9mKqDc2JcLNiQQIQk9a4uXqt0LvOt6qRmLGnCUeFzR5n8P+YWAPMjBNB3KKWxX0k
SShIwGJYNQyYZa3jTGIhzd7PMMhg109fPZk9erVL39Uh5WcGjAsZW68jW2zeqgFr
UccnNVogwkuY0wdydfIeSYzwGazaHURUe8qrg4pvXRoVCSpXt1dyvQeTDxOkq1fr
wnVPjE4hCFecWmpx1qdIDSzwiiSAaqPMBLevkrx55sKYhH049HigBJD69WHDdWi7
kdjiXMlIqRO3sDemnVfS6yv/EGy/yPemfIWRFA4x4+Kp/y163w4qt5HDrFvMaaks
Zu79KynC8TyKaSpnM6U7v3xc+G0V0y2g4d6dWDcmPDPahUpoPaQsN9kW1jRYG8ha
gOP5UScoHQlnd18xLrDHr3ThvFV3yeq6LeUSxlzt+En0PDeshDCeUJJ4XUpsC6+L
jqlG5tz1j3RLp58pQQliCSKE5UHGHzFnK9CNouVRPBV2iVrHPSycxL2y9oLmbdb2
8Osa8tfTQC/7MQ6QKJEAw5HiABTlZZQsQcwEgHsApcd55oR6SSPdM1214zLceATS
zJAUc+OABLlJWS6cxu9uh9CMOBQuYXhbXpvxcDpy6ldE9mn0Jp2o1MIq/N4oJTPU
tRBH+ZHpeNL9mVb3LcrXCB7vnKWRZeJzPZIY3HJsO3dQmz8Pr4D4TEkVOVVHcoGw
TLgvqYQj/kv/6VX0K89dCv/KpXeb0TU5DPBpqXmI5kG6y1RNJiAF1MoBHb9JWz0l
li/Es0381k3gfcYHgh7FcNXLasfHFtvB8dsqt/9pIZKS79Xe4xNGi/9VEja1XAXw
Mmdgpg3371KVWYep37tOuejVqV/uWNSXQef1Rej1Mf8tS9k6+6gbWuKL3SGh3wBh
+BKuIiqVo3spf2iTaa0ffCyg424cc999ohhi81s8MxwhXmKLW6D7XhUrHz61OLgH
+kYPTeBJFfN8gHCsylk8SwS4VMXJzSbghFLHqo+PRxhaTqBspSI8l+gIwMsQskhP
qmivvPDVpX7EQ074u6gQxxMDKcO8mTpTFq3d9a9UClHWdCAkEFjMyBn3n1fXEJue
hTTs/ll3V2cwWIrlcvLU0VEYePfvO52IJOGCYyJMmxZyusTKLe68IOPGrLIcas6j
q2pk/EWYHEX9xvKGWzH/Hy8A33a+JhWqW0/8NICHk6REbi1kbf0OyDx97PHn8a5x
dA944UgAFhH97sFl+V2u7dnlp/pQuRRTVlOwwzQdTl/sZ519ahKE2riakYtnPWfP
rTxbQFaE/ecdprs0t65SY+eF9TjUL5r89g7oGhzbZBt8maj/YdwuziU7mUrZbgIT
WXZxDwV1lCXDaHTTU3lrS86egElyX2zKPF9ElnGpf9YGLkiw3CjWpGUMIihqvNDn
jQxOnPfWpApXQcWQZZd5l4caGUT2yUXeMNpQ0NZAgrvf58Cf8ZGxmshMh1q/C4ti
ufYeQvp7jNzKCaa36vxL7cVC+utzLRixzzhDylDq/ZiE2ogTqXgV5sUflqhMCIn6
OIHyfCKIOjpm8J7Xy8clr6mpoiSjOo2hlRHzzyW0K2Tr8pvmy4bq4J2Xj6zy9v4F
Qnb3OLWLBRMihm7EHisKfNAETqKIrIv1cNkKyuxFCriQC//BuYi1jpAPkRZuI9Kd
IJ55QGWidKvNf7LYIGnyuh8r9lcQy0Qp0VW8ApV0uM0GJa13/hOkQ3q51vMFSmtZ
aIF8zlT7pIoBJKkjwV5QXfQVOpkXhgVFOK0ypH63sv18DOJ4wcPQSqjdboB8x6bx
0GP1GQjtuegzhJThwjPt97WN7ydrXo9u1wZTxCd/jdxeqq1yHrQNW0H/MIN0v8tx
5F1NKMcpzkUOrjBUJ9oiUNarV50aK1xQkluMdTIjJzxrA7aD7IVjNmjrWxL4v7FW
i8bkOOfG4VhIuPF5EjjOj3Mo/VoIwFmYggZLXi0UGxpY+rc85ULV6pEsmtxwQlOI
3BlR3gupKRJA6GSCl8U8knGQWoL3OCawodHeilSi697EgFgEKWPzxvBjRUaF3sJG
B+P9ehDeH0qncQXSusVZzHZMvwySjuRehtFgBEnEkq8suZs7m3y0mgvqupbNFeFG
Yv0JB+P13lF5vUN9efG3JNs/gmSna0hZsF4O1R4Qj8MwTse1vnSucHDAq5c7jN51
cA3jbEyCkoL1rKivDsbxGOR0dKKuMa0GPBo7Coi0BZrz+N3pfrH8IvDRI0ckJayJ
9An6cB8yp69Ez9kaZ2jzofAll/LZisuBL7Y1Vvjah61dxzlj6jPHvtKL8wHUGvwa
ewUJ5bpaADvQ1D8/z02PZSnGCewAGWoLLEWDxB/2Qe0kCVI1km1XcgBLOpuFZBaI
HMokf2QAM1YdP8ZKWLRtEYmHOrkhW9e42wFtJCn4pmy3nt4dP8JJBMthrUJ8U46J
BW5Yp9YL7+UiY5yFDVQJcvSsJRwhYti5BlQTNnLaFKrU/b6ImX3HnV+hwsHXF3mD
qytqAuDM/6BUjHNDrnpnISeh49sQyUbITCoDNDoyYdYWZc28pEET9OvGXPHC8IBz
StC2UfA5SMuBhAG1SyQ6IfsnVbW4ImNRhdV6FLn5hFB1p7JMPLHN1RHeqRGEysKx
XOYp8Fn1ygpn5bSATnrHmq02CQyy+cLUagLRkXCLQ4hvn6rgYVkkDd+SyTihwmjh
xfTXoEisJhw+LgTw1DwGr6CkHQBDrMat46YMZlAQsFsAA0y9L/8ogimiO3yB6JGR
+obdt1WUJi7vncCw0Mw0icve3D15rzH7ZxniNSbhuIvS8bA6LEqcc7pz/EkDAZe/
B+dS+vTr+4aDEyqYcqiNbjofyvPHkDLvxItzKjoUcAAydz3ZyiO2/bcI41MqChfA
jLVWB9UnOHy/5XycX9XSpm6vLY32kUcAnyI9RfE4sQAKXFqzsvxMnVQWreD07Igw
LmARveQSztuobYK3yDO7xqnxMi1LGYn3sENDcfBRYK/XvVwTPO7+owkez0O3YAw1
9+Sn4qhkEmo3UZqm+3z9ckqd+COjDT9F0DgPAtkdFXryIeq03/pV9wK+zaRMx5NO
08JpIPjIsyysGclWI+4CTDTxTr8hZnA9OG9LR3VLxjyIxYaZ8gbKCyJv02dJbXot
KMmqvp0ZoxIWcd1goxmMaIWg2cdlqAQJIVMUU5wtzDH3Qhf0cG9GMmXEyhoa/7e0
iOzAYmAMOIV92Pl68keuqnEb2g527JA2sGmLrpE7fWVBsvCx8IRox82SGdPGXRI2
YilokLIi23SrMw8PCkwxszP0HE74GAsgz/dIRXMHn932SwIiDGLk/lKPhk2pcycU
LkLQssSodvguEovZkBhYmKy7H9TZfAshtH6aexW7HL2marfq+liUiEzWmOuB89ZB
nsYzBGPrMZuFCBeYdhbmtSYNGlurj2i8N+a+zDshUu05Xg/m2paubfn2T2eIFj1f
EBSItwcTNdyeci53UyU3MfabBtmm5N846ep5sv5J9J4ipeTsA7bA4Ynkl6fQ/nUt
jEe+GIjOFb46+muiioQv1cDJ+8iLx6dvWXSM8WGiKxBoyCwE2nDgK3rAn8sj9waU
2lgBXWEeYZwtEJoj8IOMxW+yhrbBG/RmLIMJasXDWfyJXoC6GeV6IEbh9ATjGq96
3El5G2Jsd7rjoLsdaLdL3IkVOAomeRYZ2w3q3xTGhms7J0gBd5ijaL3kjHzdhkhg
N4QWlTroHO1krab2On86N38/Aa76Y9+eDCPIN2KcY1bZJKrNMOMUw+6yp+0J3rNz
VrMFd/6cuM5G4cxPI90WPzr8jvImTD4p3vdIXIStuJxjEIeSGBqsXyMtPEY/2a4U
a4X/KzWOcu73PL/TxRdp3Imy8q4/qqKfU/BG3CdOGYgSEUfI8ZmXA1cvXE45axos
nuB+FS2NqTZy6V4k2pl6dUZxC6JJ/TdNufTYg3TnpPg/lB80qpT9eOnvKKUUrNRf
m9q4oO4qQa5NLYKcy4ac8w3N4OGKv5vpNV0Y+gBEZMYMJoqPtVR4z8JtzI13W0py
fRfTF+Wz3SQJSEuYkJjKH0zeJiNokgCgGSBxQh2IG7Ho6J7rBT4IDLgrEtUmVYne
u5Y6YiPmUz6eyV/o4l5yvwkWITMEOdCwyCWxaI5qCctNuBmhaq2ChDuenx3gzDFE
gg4eKz+Ds10HShqH1mHFRDZHcpu1ymALQoUR7TeMaenxmQuHX6ocWta8i6Kq4IJt
rSKAQlm+sJTj4KAp+RH4EVDoZNWYaon3FqeghgYWYAaBxE2O9SzJh5VszBpLhzXn
7i8SQO7kAkdzcjdXD+Rq8Ud543qCCZcLcBFIiF4Uihi8J0SaJF8CrG3Somot2IbL
x/sFdLWtY0O7zsrvy30bR5KTtjaLmeD1EkU7x/J82yNQ9qBXg5mOoj8Y3g7Orwch
FwuTgkNWriIXqqtP1gpZl4FkcCp4z26YkAKgDSirKdAuQHPcP2joxsX/0jpzbe2W
vSWRRJeDvX/yIyTkf9EzbL2+Qvrn5QqDVfnVNiiYhrUAUA4AokTrr3nn7FCVxwcX
+jZQMaXQao32hmp2K+qilvlaxhMNZR1ogErDSqPclakK9dk63pwo6mBCy4lwOS5C
m7OewOxvsQriN7pqOFeswpESyT7SGQTM+YjY107a85XOTOJQ2jyMf42H4kWoZEsb
ibVAT+S80x2HYQS2i8/DR6tg0vwm1qdoIKNtXwXIu9GChQBV/dlmdGWSErlkY8Lr
5zYXFwAQj/LTOQq5S07cMAEiIvbDCHqdEUHl/GUKupTMEyPOAFQW+ZhPrXO/Qc6i
MFxLIAnebNk/8yxKZaDsqoLvUqTIm7YxdVRDSo4RYn1DVZu1f0/hwxY4zlfWHCg7
bBW8iTUK8O6vgOsQAho7Vumq3qpd0RqkWytLmIBqy8fNqmk9oGlA60hyPkSCo7xw
uK4MpMLUlAiNaacmvcTBLk/zDxf6GXaErMzZKuU4KcHEmGvjnweJ0UNgbwBYvwkv
4+T3Ln3lzCry/AJKmtSTQwYiT5Ee+cz808zIwOhFxCUwXiclkNbStv73QM8u71xT
7xpMbXpBSwzTBzn/7L+RrgizNsYkzgR1ETAs7BPzntcqRUCDB5gIOhRFLoPBeR5U
6SjUsT7tVRCwRNA+namSQvsrZ6BRdiQzuVWVQLUn8si/ZxUw7rE0+JmdBH9KZkHZ
X15l5J8j5t7iAD2xN9hzP5NH+2Qcm5HIBcOh7VgNn0z6voKLmDuGEZhYl3nPM14a
zXuqRzV+JXLnGhfXcet2R/nuu4VbZsSYn8WyiqIs/lkX3kPzR1lAC5Wtj+ckMfj9
gb/avxPues2g43JgjSnfNQeLnEqyVos0tBQW8RoUn8cDiu6wAT4PI2JxTCzE2cdJ
82XzEZST0IlPxwbRgCAG9GPFz4q6J7xZbHlgSlLGHoMOM4dNd+hYbgGspvuHOXeh
ky3oXs6FMJyx6lvxitZ1j+rC5OVELUkIjcU4RyImu3KSLqUtV264fcyBP+/UtZ9P
+cxf4YJnhDF2qXniFNj6rlVG9WNFG+842Zc7PX6j495bjlxHU0F0vc/lbzzgs61g
BmgBduS8qM7SmewYt0jHDtW/0p/QCfPiboWDJ9foYCl49pYSBOw8AVJPNKv388Is
msMaWMZ1W8SEwUtB7CZQv6LMdHqrq5XER4Jhvq7ChGWwxIgEyGLRvugZSFt2Pwis
UgEJqnvxKesmLYdqAWEuZc4bcpS3LfCZxnY0rquxnHqPKuZWg2X4bc1F/moELSxf
12qtKwY/eSpWZ2ggIkltIWVL1fEHDpAnX6MReaacf5Ql0isyoHV97TpCgscovP4a
woYU1fiSsmRkrOfuuDxmqPgthKMCTb0MS+NOKU7Ggnva4HFlDRFO3w2Q+NOyKvdC
C0/YBF5Q1dMFDg1c8pa3gABk531hjjIH2uOIn+A/oG8puVfMt1fW6P+39YfPoSI4
4Ajgd3uM7agS+f9HLdkMacM4zxE7ouAineixmDtdG7lhL0Askl4YyypZ7/wzzS4k
HUp2QrrVjqrOQU3SQEHvYDUhrxpK2XoJ5VnyUaz/YkqymtNkiPiG0meO8+s846ty
G/G7KcCGS2PczqUFFYat3qmjuxTj8HdMcRXD4I8iMRDZ/IlZPBZKowoV6DKi4FD2
s/1pm2rm3QIPldVB4hJSWae3LRJBEpdQw4MIX0t2nyxhVOGbJAA3wEdsp5voRCVA
mAUGGgklWNRMZk7Un6gkVrBmPSGGto0aJ+mD16E/MMr58FfWu1ziHKj6e+hFGH83
DJzGgtIdWs4Zg8JO/r3a/aEPDlYibbHg9I2/3Jn6q8NULDGgV9dgjyV2+SaHCFRX
X5aGm6v/Z/FNVzGmEXanYwNxkn2F26sPPvDLm6Mlk/GPwhQMMA6S93jyj89+GlNG
Gcr8g+1qxIbDQ/K2pZAQWTKzaLkoWd1t7t8UbdgT7epr2HtfdYdylgPWsk/krpat
RlO0qXX+rFtsYTaA7YuL84MM4SUI5mWSeiSjxycTfFQKo7Yx91dEmEo+Jf/ePfeg
o8FIvTenS48K3pbl6dIvw95M9zos91U4hWJ+pMKm03OWaq2eJSsKcUDiKbEyd5ie
vjQ9vEcHr7ncDJ9xwym3EOyc9vJoxlrmSs1V4/49reIlvrLZZbiTM56ODZBluBLP
+0lOHaU7xPnt2wWZWkpGT2ZNcsliSitMk7tEpX2Lew/al+QGDseaKuAbk1uLxawU
Vd9Gr7tkoGUxCv6JV1XOKkPwtrNjViJ88jvkMlJs/9k2xfZ+c0vL44Y1gO514od3
4BK9qKdrxM6YfoWJSciA7/80E8yAVWtqQzmWdxkDq7xZFaZgpWz94X8DT6xzwcBM
ckqErj43lPT9Pp8wWSiiIa+2gtf78+qoR6JZX1H+n9C0ST0bjvYaT7XW29IW6YGR
6iCvh/y+yAz7CzLc1efnqVT50/lh8NWL9zxKmxILmUritRIidC5kRGaCZzFf8dtO
9cFMq2bSj8aXgSnVvU44jTwq6cB6uhDNF9KtVJDS/Aa3mPVXs5H3VG3ZF7ucJz1n
MwcCPaLCW6mSkto+atW7UEB0qaikP/H9kE1ArOCjjJVRAlminEU/Yn9YtYX28UZv
suj4KllQ5BE66iuZsicBU5V2OpZfoENVUxP3flpl+NkDmtqJqM8isouHjtQprlS1
PBxFE1FGGemwnRZEzjfU2R5xT2JBLH8RKJkkrPxMoJ+/ee6P/j1MS0Z4JaOSgLA2
Qg2Rz+XRYFysEFLNxYfcutP2PF4uTcwZTEK9OsCEOwLcxb9yPgJQeksRVUqIsF9i
AiUyP9s4Iyu+F4CGA0cKVg+Tl9yDrUtmJMyfQvQyH6qX0VCWDVkO4FwbNtzFNhkG
x54/2mGF8eOqAhO/+EcY0DZYOPVds7/AnxXM/occJI0/0sCdiOZ60D+DF3DVgeKe
3Y+JDDcEKMuQo29iJwfs3a1SmdBTM8IApdViNDCP+Cze/ozVX0WXkgCAzEXnaa2w
T/fsyiM64ItEwT1aH/8+t7pFfrOmq7DHdoWPc7dqx9Iw0kd3vnXmSLoAgyRDBEAk
m1MMWII87Bwm1Vb0e6f0u3aXTtEkIRqTa7eoKhkaom3P00m84fnqJXG7cKztqv6u
p3GUpb5zmdXBs/CzDlqfycxNFatButq6wzPcTaZ1kWQPHPSOehza+33LvAi5b23e
b8aw2yrimJ2pz3CMpz1S8T4wZCspITlo4pkFzTyWVH2251LXxDAkpMB8DK6W+cNN
o7I0oeFKzcsINCAsNmlSr7qNgmwm8X2IxPm7W5XWVj0jHdPZ00SP3CpovSZyG/f3
JFKIKRqEudMCkR/tmPMbH6EA1bSda8HcLap3vTjX6nx5imuu5rjHbyFrabHYNvV5
IhUOaoNjH0QCmSSxk9N9WRk7d3TczNKKdpYp2RHQjvTjJ+hsT3YDQyi+DtsCrc/1
XdKM+SAD0JwQbkGcgK2yEes3fkH3kWw3XkqEU1jIwxutj8csO9IE1Q3t/+0Ilg/h
EFu54q7aEMqGffw3/F4lOsyhANJkL2/wXTPtKhCI/5ue3VI0rAKKp9kYLlKf5ZkY
omsdoQEqYOIYyPWrPK+U9kCzak7+EINrD5/J+LcAfimBXiKJaKG6LU5Z9zrvjbBv
Fz3ePd0TaxTYT9INhJKA06gIsc1vINoE0Pd7u1TZK27pyWQ5KzzoQvw8HsCpQUBx
a+x8C0SzrWt1aUIHqR21FjzvgDVGxvFMdXfZ8IQ6Kri2DDpMufZLOQRmYUfRmNIg
1GWrX4GPHOSs8aSFrumSS/A+KV5xHmj2uuY1qwsKU/JUMzZ6BKeQb2MKnKsWwR2U
SsLdtzGaLpp2G9DPCgt86ZjkRvOhDgmrEvcRb3fdEOrz2FFMZWz4EQDCAU4WjdgI
Ztp3k0/AMiKLaBf1DNmSqA69zADuwolkdD+Lr0aArI8S3xHLl2Lov7YOrwXTbuKh
UQLAorcU71qfmP8CLD/gunf6jfWJEQqNDZ0Pi/F4ndiFU7XpDtMQntswJV1g1Ula
AabGYWxCANNEvng0sIj8oCdtf3raLotZZ5yyKKJzh68tYtd3kz/U+zZo5scqGrNP
1YmbkL9ne5k4NUaZXKZXE/y5BDmRAJy8WIwlsoqQSlXTWlfUyl6cncuDzGKuZVgM
8p1737tugoqoY7CP619DwE1xps448r88CeyxmvjOXbAvMcYYMDaQUEFDaMvB4jr3
eqnDDQyOeu2bEMqlKuoDONw6Pcel0RazZscj3M+0JEpH8CXDAKh9cJyzHQYZLamw
UxjCijtp7XF1UKpgdMwwJUMUDcZmpWBgsXFkLN+Etn/GPPFkynT0yHoCev+y1rKj
6a081Z96EKlVa0Q0itJo/oyGZ4EbAt4DEUhzf4IPw5Nqjq2KGrLfqPa3tOpPBy+w
7gGi72WVvmlbv3vdC6Jn1PRRP9QPS3Fs/ThNUwLBF0CxrBMMCoBlTnusZM57BZup
vTxs8mIgGHezfhzYvpTVLHieJUjkwjc1zmcs9og35u9/5b5adXVyfuuC6svcY2nP
VM8m/jsrC97Bt00grO4GOpRZHfDkKTINbxvUCHPVW7bYpK4xLMkzgYif2kXEgReq
WWQG6E2SXo9h5RsYibuEtSDC2Y4/NsK5BpPlCTtth3aPdGlK58Ix8t5sUH9qFR5p
M5B9GPFtDPpmjGdhUKRFk3cvC5cOZ1pOG945uNw8oSKvM3l1IuPVzWLSu3OQqfdt
oI931wntOzlw8PA1ywoNty9nbbOV0OOg2ca/8SpllnAXHGtW9b1eOCNQYm8IOvMc
UCk/yS8688QkSERFtYoZ1UhhVy6ydwNUPHWeTGVfG/sES21ORfy1qZWO/Q70kxz6
Rso1Cz4Ex4jXFqVtvdlvk43WZhYapb0jgqX8n5Z4f3mB2mFVUdZ4lI6iaj4hJkkw
rSJWmraOZ3ebw3w29Rm7WOiPbAqsiVj6ESKJ3wF4qDEIz8Tymf8OP80iPWXTyA1o
H4JozBKKnM0e/5uw3chBv82jQz8oT7I22sR94DuVjfglfk9wljBKnhP1JP0eWbzf
TV4DCNaEX75clpQq+jQbux89qUs0ofrb1eY9Gy8nIKLsMbHHa2zEFROZnSqeQy1i
Vj2ygCI259DIlzj3IZFzvRdvrebNVtLYpljX4EhfvCyhrrDGX+K6goSD7wS1bWyd
yLhTFed4YAybWBa7pSRY0TITnsBV5EXdIqTByhs/Pg7a5UpoV0L81v7QgMUKkfa5
xO8p9JmOTq0LU1KzhVbbWNiNxinrK8K9XRzASCO/LHj7TPcnkVq0L1m7Kxw7MniO
vu2iXOFzUEzTTPSlgh+98l17HdQcmXnTdnvRQyw/u8y/+YpXtDg1NB5b636MJ9mm
KS1GIDOwg5YjaXP6Kb20eDjWSa6T0RkTdrRa89xx5J+gMNr4rgH4vAQIowx8+L3X
djv8pbvV4YcRjKzR+ZaFwXEMyUrm6UKKartqIyS6w3RND3SbnMNrQOmwhVyEn38t
Vdq6r/h6yNOGzIaGLVVz1qn8oXpPmvr+uKeR7h7Gohycn/tFdyqsPLAc7fHWIDGr
Gh7BblPf43Nzi7Gc3+6XZH1XfilikMYKWQlf+aCCqyFEYq6xQrjsjonWB3XO9RRw
f5Ex9jHfuMQILKvI7ss7kKvtwMqf8NhFFVc7DIrWLOAsOSHaaMUadlLMVG30oWsF
1Sca4iEnNZ6qxU+lhd+dBP7KZgGDYQdrCxD251sqbzMKAOjvgGr2OD8svgq5+/YN
tcpBnAT+6NZ5v5AVnTBMDNi+9yKBkMEfPnGijFwDZ7kFP0oPNwZNaaSSsvxZcdSi
qAwiPXW4N4YH9mD3eHefFw1WnAommERNgWTUUv39PDWMZu9qS6ONi9lpxCUB9dGQ
1zteyyYPduijlJ9mMj2JyIbRZe51uxSBO5ROd/j+yzwT7kRuNDEh103pd9Cnu/cw
rH6VOh5R7rd/yhnEl7Fmnfacv2wNZYATgPt+Pd/UXUWMSmw2FU+Hs9W/0JfGJktj
99+9OnFnCDvB/qX9BVwbrtYicpYlALlSU6pDFWGW6gGPua2BvZ4F1ly7i8T770QG
pHRerXoIcdotvLJFzD9CiGXw6HRAPTLrgAXKwAKdhrO+WY5thjbB+N2NsFv14Upm
lXlyB+If6xg/iLN7yUMSw5hmaZxsz7R2fzRZhm1bd9mWrbWsMIXfgTHBoqqQslKu
6caKi3E6Q2UTbGUpkr9TuaenHFmFhk8nIyfm59cQHHL9yGGpF7eZP9C5/TdR9EAr
YxTJUVttOQ3EMGaKkjiDwKyJ3UkC5cCw0jr5I7R8R3EbRQhVLpU2wWVZn1yzdwtM
kC/yGPCh6wDjvkQpsYD2LzdUtOu3v+G9YeBpOwEUw3tfxLlBB2nowX59JaTUfsq3
P8Lx6sG3CYau7EXUFr2sBKowD5ZJNIAi98TcysJEgY8rM8KsylRXsmnjowOQJOcA
Y3st1ps2MueW97jpmlR1+cU8ekRXIU+AzF/6KVrm5T/X98sdv+xyc5/ytz55QT+o
S9xGD/deeE0OwoPv+oTcFgKxBMJBgB+T7rxd4tt1oRElt/JbjZKQcnXAU+CxRn33
gQ4iaQ0h1z2n7LO5rlpY0WmRm2O53XuorKL4/6X0XC1xvj1Abtva1xw30INTJyq+
owLO4rJNmCJtnEd+AG04Q5T9QZdJaaDG0KUZV2ljL0kQNg17LyT6mT+TYGt9m/qP
37Yx+3nzr06lz3Ojrgu8SGnmleVei17nNqt2yKD26YD5YuLkk16p4snMC/T+aN7y
v4voSjVj9Gk/ivrPvRfSu9R7raGBqKyjoxCWaX/ZYwQyr9vkfB/Xg/vrsWRk1O85
TRGgYfgLh88T1dikq7VlxMMmkN/6xRBO4hGb5MxqkgdtQRJBcQRlc1JRp5XMIMW2
NsvUvSjpJ03Yawkoj2BX1lXB148UheTNa/HBn+8pHT6BYssezutzZ99rfule3BKF
U8XFq0U843kXZ2WfgurGOa0w7nahdZo2/VTtBYcJ11eUKsj9/A5S+1WESOgOE8uy
QqeDcL0VGwFmLWtAiq1Ky8NwdKS8R+Wc/BqaVxFcUCkVa9cYf7zt99yZ6r5XKf13
rA1VVgNYBSbFu5BmM5g+00WjNjuZyD+JBQP5ODKjm0zzNAKqxlkGaO/SbZZsoJ/j
Pe+tEv5BfP+ACCLZASXexwxtHq7OTfH5Hq5Ke36EjzrcA8O+jpqtlJ1kfo2QyXG/
Q0SXFTbaFN9mrBpu2qTm3BGNHx+BiWAXVia5tK3BAG2i9rXPMlZQ9O9HdnpkKf8V
onWUcB+KrZtZyRjYV3sDcvl/GCJdJgeJB57mE87nMEKXuVc+1Wc7gR+bzCRpohXb
WoZnOedIFtMVgKn7Bo1kGrAVedXF6oH7E0eHCwKuyex2lSyZVI3UHMfSIfTkw9SP
WB0mbIFCxELbkDuZbk0A4P2+g56QG4qVNK8olrH5zLTAm+XVygpu5Nv3GaX3dXBk
R8vweB7o0sSiPWz59+D9hdfVKsbIL6bGuJPa/Td6rUfYGWh6+ZGkwHgjYqcpBYgP
bFwDiuYfvVm9zyddKKptGBQmpVxr9vqrFzBz/r82oGPlwbh1lDnOuEOWIuztNXsT
Vc33a4fjqZtqPBOdro5ksnvLvnDQEEfDToyJxCHuGtfRbggqgJ3hIEc9EUrFsk1+
FSN0oDyi1kLXbiDlllY0lyn0HmEsO67Y2UrJXUwi4wBF52FiVN037gYp2qBnciDc
m5NuoQdWezymZD7JENh/zExSU1jWt7fiRy46b9stl8ie0QceOrsth23jY4L3aO/8
xxvbWtbAzbSBu+8AVWdklu4al0AgG4yppmRO4Sdp2rnxLAbkRNa0kr5X5tp5EGY/
uceAhZ2dvvzyQBiMba1qVulUWeDFb4DplB5Qy+eT8iNwH7bIHyc5U0gce5yADZrR
vl2iW55LKDg770yAR+4uOmOXJBfsf6wTvXbyqFaTmJFDOcluSEIEaf56kc83scNW
L3x6b11kKl7PJK6RnbbDJWVFE026We1xnblcmu72BAV1ljOB7Gd4c7qYORGEndg7
e4CDkMzCtriCW0h1fNGAAEIQr1ARDsF+PXEJoxvVmuXgXq+kNcIPCnqxa+428PCa
hT2OreL+M6+bn3kYrS9VAPobQ0BgZB0RbG3WsnR6J3WBo5K/I3+9tmuUL9v//0eF
VAcWy5jxKxcvyZUaGmILTzSuAWyay7VBvx9ZLzNvCPFaqUjV2VVS5zvzf6b/MXKM
Z90h2cH6ODrw2VpxszZJrxaekxx9deO3VIEyVhIOf91zbBBGAUwnOXuUGzQMQ5mB
l/NP34Ke2Iq8uRKq2uMqhcD9wWV0FS/NdZQadgefCjYt8D19et/zwSHalUjMzwTx
eAsGoG5DHjS8ii+ND3qNnQ/Vuk86vqzBBmIoeGGEkYX06TdKWtvJbYhEwSVV8EU2
T8D6c7beEComKyQud8Mnqe806fbE/KQ4IlBKPLWA9gUH/oWUWZZlrR4qykJk2P+I
22QfjlntzuFvNArI8wpzw64VBG/UjOX8i8Ywsk81/FZ18L287T2FmnOT6VoJy6xb
W3d39SoPPclk7Jn1CmhaCxGU/3LJUPx+WhL0TV866MyA9YubOOhuUwbpg8nM6FOk
QMRIY2cFPw2i/LXCV/zMFdQlm1fmyvv4AnOD1uksCfDfy0WSYsKomcnnwiqZDuuy
HKarwp6MCHg836QwBa95oWy4lnu0hDf+XOgO3zLDJFuqYIjUq4t6+BtQlN5K0l8v
brMQ+YBSAtusu/s5dCyameGJNW+QppuGdnu2GQYKGWisTTnac6i2PsHBM2LOnyUk
y2PtrikaflQpZveNbFqGw8FIvh2u6kBKpF59epfhiS6o9I5V3tpvcR3MkTF+B9pM
weeUF7npOrD+BOH6GpJqezN80narkx3AbKZQ60YMdw8TLW42tqCPr6RH930wAMoW
XB+O9ggCO70F2Vamt0FDmOXswrrAGgYy7SAl+HFAfsOayZXH0/HUNZHAcCfxVn3L
xJhKdpVqaBLzQj3eBaJ1kugY6ltH637U1n/Upk7QpkOGzx09YbfSwwCObQLqpvP9
lOA0aWXjz3HOmnocqGPAjJjLHsCt6WpF57ud8OsVe8DfmxUsppTUYKfrN/MjhnLC
Q3Vg4+3COn7RGovZcsAEZ1RmuEcF65TRvFEo9Ok6SF2n0b3gpQlYb6EZti8wQmSv
n6Kdr2mkYGMgLK9gcLJBITVfwkbMF9PEjw15B8arx9SbZAKUkExqA3ijBoEbgq+H
AF/v/DCJUIW14D+2bAgIbjuVzmIQCLhCP3u3hQSR0dOaSftIy6Wd+aKnggBI3Ui1
NrwNYylK4/JqaxX8kebie3ZCbbgwjINf23SZ6AgSwXe7sl30GHnZlmBSs1fatf4w
9/5htbCpguSR25QqVNTTQF++ee+uLpyjMtcmNunBNLZVOfpeZAigkZUSE/N9Q80b
z+qyTS/pn0iDbOil00tbzvQmS5CuxJOlbrULIFVRPALsMe4Qv1LFQAHBjEGImadT
Z0SzTJvWki3K0t8KWsw3J+nEyPilfWaOXbIVUQo3dvTDot8uwhjJI9HSner6gDJ5
nVjcL4vS5/bc+yCCkz5eHJrsId7XFNoCO46GUPLL0OreiYVwYRh7KAAjTVRVNavT
O+HQ44pWTRj6Q/MbKcUy1mq93IYm14TqEUrAw/OfM47K34SFURKPcWeYyAhnccyq
rRHaZhiSNvlVukb+0DpC7S5sSkM5sMmkxEyIop3orfWoCQaeITFAiaTsyweX7u/1
Y+W8GAocT+QVYNE03XD3ihza/TZK8iEb2XZyCcDGubmDBTzaS1DOFGXXugHLss0J
bOkbLqnHvT0f4Tc1sb120YLsXdh45Ew3/MKb3KHS7f2xdFlBbaKtNbU2lxb5GBNU
K13nvZaEYeZqBTJefOOSN74xpUF6cujBA5mjL0DByBV6UjmXPYxBqaz1PiPLD6AP
6JovqHxfXST4j1gBSxmI9Adm9k/QdzffWFng0cvbrKOb/qdbwcwWe4YKpvS1Pgry
TcL3kwczxKAB66imXpA55+Z1FN5Q74AZ3H1jQ9LUdUvHCVtdNz61S8raWWanIBAA
0/VSrYw4DTvc5CSLWhkM6q4dF/SIGf4IuAO1jpBEgKVMrjN1YxPivxg7HK5wTD7Z
jkcjWLmPVVVve399/5YlHl57tzMR4WiGFEIBRewLJLpQwrAkFM2+xz7acNbg4n11
n7aOZ9C1HQ8dine5SQcSbgPOwBBKt/k6v7IqrNKCqAKlZWPs197fhHPJwhAd15Qg
pAgwEW4SlP7Zfd9sMzjHSD1tj9wxTKASd/tTTuHnSp4YL6Pf7CEDRl0LKc5E9O1h
wXs3rRYADPozQnls3ToTalF1BjmF4o2F7TfLfKfR963d8RMNMneQDWgFuL5VCFb1
S1jzcfnovsUpICz50y9V09fFppz5/tPjiJenA7Wz1xyKPq6AdFMvjDQv07urEgn4
bKn00binWgTHoNkNTYh2IEYwcYOH2PWogGzbvbZA0d/NKoBHGrTvR6wsOrfoXAZP
XzagORwx94yOkyDYHiThofIWYuazKeHpa+vZ89ZQL0Xkr6b2QOlRxlhlnENwc9FS
KFP1djRwK/vvT7XYhWIj4ulB4wSkpgUleTNYSzHyolYfDC9wqn+QMysbfs3+rU8f
+xVf8auOU2FndzF2sNaDYcOvDKc/F8yBpgoJMi6u01HWxpYrSO0R5Xl63taw4SO8
LJe79Pb9XpJdaWfPu/vVoZ2RDOZlD+/+wSSbHyhPS+dBKwvDBIMy/EIFA/mTMLFI
TWr4L2GRnm/4WL6V/bNSD+1PuXcNXj281n8hEux/P06vagdXiB/DkS380OjAG5ER
OBRklrw+E8OzVNP9Dac+EiE+y5CDxZU6tn5/xJh8HGrYfhn0BUgbwVHa5ywIpt8Q
Nf45UamcDBrY51BIE1VW9clgyQqdTIjk7B3pXlNOZeg+Dm8CHIRhLG4wzeD3R2Np
P75rk9NA0VRYu0WTq1wd5qQZp3MRli0f8L9b3K9n9Ov7yoZpdGtGfZvlcV1ul4wr
FknN8Z85iivVDHUGPNUY8+FJW6TDPIOBBNSwBosNYy9YhEMiYhe9ixsM5pBF3E4b
rScqloHwoCG9nMGhh19fepRBuo1cYEW8yPHeSMqsZ/Gu4FSOw5Khtnq8laYNFp6J
Zmhgq6Y6ZOwx0nOxjVA+rmU22TZzKpUiuDOJAIzBQ/aTgl2vfNRZ8dM1kCAhDjXH
ztzfgA4k7N9x948D2eSMOep7wZzBITXpvQ4zWP5Bny7R6V+S0my8COmy5yhEyeJs
D/gkOXP9TenCIdd5DzYihhQdOrsWW1EoRvP00Zq70aE7Ifnt/C6nHarSSiiQw8qp
bxTBwztpv0hAyj7CXe37ezRDGb6APdFmJVPDabGZZMrsbAWPJXRo7RFn1cNt7LkY
/16rrpyNLeGyntTDdej5nuumm6pVBQmQ0/7UXod3503K3q5kFGSD7U56CD83cPHu
X2uQjRF/ra348vLtuJlg0r0QS/kQW/WpGq3Nx9dRGdmlWltlgwUG3KYVYqHDi9/1
P/e8Xb/hVbEG1yQXEfQbCrt/mKGMJsj/xDDxE9lmu3d70WTS/rAYFb+cqQdFOXtS
S2OYssDDoB5Ololp/YCdyuMzIhD7dtp9VM2HXImPe2nMKXyav6XA+ImDuWR525GK
9BVZUJ9PJAtNixBAnsTZ7u+Tj9UPfBkUDZoLDzmXTwMUi5tD7DCOQ4pK48UJ/e5p
ZGIRDfDWTeIWTVTt0Q2JpQcFjiF9PHRcsOhRL7DILP+x7p01ps9QYlrgBf8dp3/L
NOyah77HQYKnjy41onPOBPp4SqsnHckSYJcakh+7W6/8BZmxMef4yWWERA3+7N+N
XAAXXCwLji4EGQkOqOMlW+qpECGl9pE76UGLNMFOYmorh4+hx8u3VCIY+JqEQH0D
kRehqZ1zWgeyvbJOONbuOOxyk30BIHvhgTsfsgR8T7kShqS+3K46dshJqhzv9pQU
Hv3Ad6VpVcDd/rusDt4V4BkyiVIZsJVwBE+VgQf6tpaZQudDFVJ64xUK47Aso1AH
UDr/BUlFqGfGzN7VCITd2cIKlLe5CkGA5KfgEovBI1KnRgch+wdr7oD5kQwMzmxW
vrRcQEPEZlpsSQMM1fFqFV7FVYOxcS6g/DXoddXGwOdsO9IyS+O3VPPgWVcQIvIo
uWsFu0MbeR/HbB1Gdx5XyGQcMA3LJz898Q0r2kVAct2XliaPsCVOryX4IoOXF2if
5BmmcNjUXStJ58zzVIF2aoxuxha6mCynLGvz2X7uDLinihA0Js44AAGxnjlH0DZp
A9dCFIwkeHsS1REFoUGsPc6FcnQjYvqm9Bu77/seXWWPFJYrZDQDuOVSMeDAHIMi
smd3AOW+1YfqQQkYateROtGAi1VV/X7BDVwbycczNWtguxoW68E/0nFp76PErAeG
ADfH1sRV6Dxzd7d5SegMy6OAuExg3IsvL4iWTmqJju2I/vLSANbyOLyXEw8qcz0j
bWNMCu+xIK7kv4uT1IS93h6FgmI17OcbYLZrhQNgYz9ZHy5hXojpBEhxNR6nzKQc
OsD9XWpqyO1nHQkDWlcnUB/3BQAn3Kg2NlLAU9dj1p30BQdEA6/ZvZN2ygtOp82D
urIaszlNNqWGm3T6JYyVBVT3Z2TLDdaXZ7ojJ/rL5/vIffNTqtPTIqBKDnZW5UgW
TUgvqOeF1/uBKog6hNvQhIahGNd3wUMIGyY+nLSfPf0jc2zsXP4irHSrWM0xB9QD
YQBwiUvdqxywdrMhejAOiCgd3Cgld6lWVxbqQOL2NGISQQN87GvI02nhANGhOlN8
Wde5txOFnSkzDoG9Uc4zLd99l5FJUIYK3otbAc6MBx/34OURcPAeA3hdyTWIu9z6
134fEyvn9GU9yy5b3W5J9sx1inv5O1oaOGxJSNqfThvWZ2kDZnnuqNthBWRb0CSl
jMlGHS2dpiAy5vBcL8dEgBR6d9BXX7dWrMiJ49IWhDDI4IKlaPt7nz6kq/oUfRBQ
DciyvVHVd/FyF4rBHdfKSFkU30hQBFcrttPiIRJcpW1ysyfL+IQaTFqLS2+Jc4xq
zR0jaibNgaIcJg7azDwQNZzkInRjNVBn5zExu/qDCfpPgGc/MfAJxPVrD4mi8EaN
FK7qw/N7JO3lmSfQb+Lfca98JTIcH2ogoo8YsiJHcWOKmcFd7/ax0ku3Fn6Xk4e1
Yj2q5ayAwm0mJ0dr6twTMAv6Z/OFvEnocvTWYdW5R/OfoXXMca3oLiijDmnDviLn
IwLYl2OYT1Bsv/haPttPAe5Iv6hanXpyZKN9UCmy3yv7LML+BbV4Mw7rpXvSpvaz
2qhlvLorjoo5SrWJfoLXsV8PH5KtflBMT0DxTTQp9VWD9eDO6Sc5ctMKwNqh+59/
ux7ZyuYy4x3VTJdPnXzq8cNaX3A49NSYZ3Zw2LedrLUvHGqxeOY2mXx9ZHn32LKR
WUxht5fwattvcQckJZDwmqA5EN/7VtywAFpTWpjP3dwrNQXa1CKueQxsc4TNHpDW
aUp2hdbSDZuu4BWN2iGLbmy8ywCLsGlFU1OPzBYjHTVuzk6UZi3SswNf7ibmjO1/
I6T78JjA1DHW7Y2jlrhtz7zvMk1gSGNnb/POHm2lb7ie09V/MOoZFs+rKH50be1p
xqhYooZsZi7NDpdF93ZoRiqfy8/gWuTUGUBPqmKIJwOW8B5WwFsrpyrXIyELUUdw
71q/HdhGie/Aig2BUkJ+GfeQtkAg7gPobFs8d99ttBE4Div2OLTZIc0DJBO5Oo6o
lGelToJVDrY+xayp5HuI3mSk4bdtYDY4Qx9TMufvZ3IZn7xnDRc8eZwcwnCBLnoH
pH7OM6LBsxrnyM6SnwcQ4M1YXrF9zBCHk3VckZmB41sgiExjVP/GFK6NkpMUsgsY
UwMa5X1FJlszAXeQTYauc32R9z7l+sZeKJU39IBVpviL+2ODfHxGYDLQieWvCUEw
slLmQnDxG2HtAtpXizUCbIBR2jVLMeSsNkpEDp5prAeTnyJGOWbs7d5+kloKU5zv
UBG3z5DlCebRXeqLTQ8aijeAyK27WIm2hJEzO2ZchwZYF2izWux1SSI0FQ5qYBpx
U4w//wVGM4URHk38Y90dqQMj2ZaiqhEhbctsLQHNiGHcoeJH96K5tj41RQ5B7wMr
IYNqDPvrhRZrxW29iuyAUDnFbaxfP24oUNfh+tl1zjU6+DWQQgzggZp13m+KwCdm
yyW8JnaroA0rpve85xE488r/JDZ6C2QlzLjqOMR1yQ9HJ6U4vpzJei0i1m5zuzw1
gJRhas+zqwV08RAsOf63vMHm8TJBSAgnvfA3iI0mSQPOELTjt4IdEqVQ7b67FGIh
mzd8C/imsqhWbQ9BnElV3c6lPZ69K853Rxe95usQ16s0mDkQbCD39GVTwiJ4z3u0
J1cNyAVzBvK3THI7vuiLI8XZw55FQmbwi5oJoz35IYxuBjuzi4pbkGdlY1VIBFSM
NAQ2pP6YoA/VW2OIdbM63SQEboXF1Q2i0y63PuYUdQBROO7WHALhijUCT9eVKcYZ
f9vBCmdfDNjEwl90iNYMJoSo98zi4DvpcL4EI99Xb7jYfhgJEAEoRzwJyJIL+MBX
tfCwKUTTH6nyJIdeNICj9DOJzxEXebsfqd+l9TN5GhgYf5dkaS3crZb1lhUea+P5
Mm0BCp9aGGhJvNlhxlgF0nrkVuEQhfsRckT0Ru4+BhvfEY4m3qTfZW7Y7us1mW5u
GvP/VLWAXwDC5KD005+weDXW5VTerjHEOez6IAtLGr5UEf5lCt/VrKr6Ir9EEuPa
wsBeOWe/WKlV0uRAxeWhFn457W/i6jjBeU9YI8K6s45xZOmPmbH6aqGzWTzuZbsx
UjdWgJXTKGtTrBqdjeTaPRMh7jDbICgKrDPoc6uhjPtOR8unDCnLzOeSBmd+sKmU
4r62wqX5ov8BFUkfrBEW6z+qxG3b7QqedgX76xROBhfEm5aI0lt36YZdT/dkR5/y
B85fjZoNYOVjYFo8m1YqXmLwFb2YTP9U+tEvj3uplZUUjfWzW+hYreslAlUj/4ty
B+FUSbofJx7bTNQkTBh22QQVxmjZVi89UPYXnVrG7bDCshI79+6wzaVmrefXSSgR
az6wFUvLYE7827ES+wEXmNhCntdBODdF5JVtQyXe4M+Ub85PugkQGd98DnFAMLpH
f+BatMDefgg0p60Ew7srrhlbP602viIrI2Q9x0n3o+1sewDE6bje1CzTUA2wOeDX
dJNaBomszj4h4a/QF5Et3X7KmziPd/65IibMAn4t2XpmxayU2KR3KrZ29Ytqoysb
fBGfUL2zDSX93nft+YNJDjCubvH2IaKttpGuzEcMbCTKP5vwAHJdWPQ78bfnYBfp
gK+6iGn+U30fIFHBEWFwqOb5P7/DizbZI15n8rLnpHL8ma38CznWzkQS05UDU9+p
a6E5NDncOQpWcLzXulYf706YtSdjASiBKKpt+kj7nPYE+LGXAS1DzZAHlEwcLEcT
bBqd6zxvJ9cakLVl06EsAP/7USfvDO73PJvVh5zWDzNzWf8NqCPoC6AEPAWHMfJz
Jt8Xuj2Alm+UcFkpaDEN7S3jhAoRNoEJzowTcWfmQsbKdcuW9E7UtGz9T/23kyiu
R8NyytFsyH+NHMJjVnJpXM+Ps5J9xsL65kK5aEsfUA7kSZ+wQYbJ/p5r+k9SEBrG
n2EOrQy0A5ZYWdEGoLz9stMvll8k0xQ/8hqIhLqTLPlPL5jEDzOA6u43Z7Qi8E0G
sOGwahXKjwlrSbTk1hLZnedwz1bk8RPB74F8KoRNV4CPHlSyXeDE3fdzkeR2DnEX
QrYp7ynsgSmIhU10YaV+sdHWc5l5jZJmDaDr9X6UtAs2fUmBVHDTXEsu23iFVgfc
T8fmD2njUyhJ6gqDduOmq4Fnmq6jLLl8gICnD3k2mMdO+2550uy4BTUR+cVx82MT
prg9kNsM8bRZyL+qbcuwexV+zpP5sNiRUFGtuz1XAut1vrcf4+sPkAXl8K4CMCxG
1y18ajrdAmqUmjGie5tErIK+JZTM1ea8GfKAi0NsH20xv+ImExuRTVtoemXZTRzv
oTZsaWzsfZLyuwC2fzRxGMjmBHyBYExebCJa0zJ6IXejp6tKLV65JTP8FX6ZlwSo
u8uZWnfPJhiRhdIDdCMNTHgUN2Zv4ofnzd0yGrrTv8sEwKJcp8EWnwof29TfLSB7
Vq2qJ1MLIrTPSZkIFsunWYSddK00kDxula2Qehj5CD56bIT2qAh8O22q9Oc/Lkhx
wHdfqz0zv11q6gkjqhWrauugjxTSkwsvUKQdmJhd6tnV/8RnB4VGIrIrRA3rS3rS
sPyf3W1uHqZF/B/Kag428j3S0/ch/QIWgxvIOtRRW/2jSyY7/DT6trtuK5jyQvIb
+hgcuFdFzVCjS1vHBlMW36yVKBu2DQC8h7xwSNZKAF5VlyeKHKES557YLmHU23Bg
k6LAjRi7hSEp0j1laCCn8GJikCfZXwSNcxrn0RDO+tTDS81uW1I8P21khgrcYpMT
oR0u1fFMJ2Ek+xTDHyoZUWDMrmG1hx1gkTX9ejtzcSSdssF5GEoGMnb9SAyndH4E
OmkMp3D/OjT8CVmJh9B3r8g0zwoR1pt4irpOuAE7uwfGf0F1lmD8L7TjnJG+lmjq
leGMwjdM4gIOvYvv3ud0s+R0lZ4Ce+M5LjzSAcnFruq+rYdeLkyWW0Z2YVuAF4/5
N6BAuodNMDQMzSz3Lr50MOmK+Nk+OIsTgY+wQareMDzf/PShdf5i5KidFIYxkrkX
nNmS3LeKD/EMCT4klW5nExCTlf4Nt4N1Pen5Tq+kPwg28soNy7ofVVW3g1KbvHnX
GIxScG66sOdnbiDnPsQlcRSt/6xsibBCPDKNx3ngBDNgl7q2JlhiCmD2MqFu5HYD
jrloEE+pESAEnHgfq4UViXn12xWjGTCzTd5ODM+Uy0OBX1Gd+eXaW/r1dQpYAIxi
0/x/7tjgHj07NBtQ/92pk3XH/xFwzahP7IMP5gu9Y0Te/npTaTW48ebuI9jXdaUH
ys5UvVxrVBp+EZvjcff81DAXs1RrrisAJnLgiwLK2wEZvvsb32rh4gYdX6ocgUAZ
faQVDS+J5OBvR9T0nUeBj61kNhL/6ztzp9weg5q9rBf3fY1d0CawHavxZQukOubS
zvua3TIDUSEbpUj/oMtVUA58Nf6RAdIzKLA7WpwIjTCgJp0DM8yZ1aEGq/z2QxTL
Tr8HvkNvrK2AXqyw5VrMHPOFcnyYLU1G2bFYd7CuffvP7hVP6pHhMWSMfwpFDCfr
H3DW/zhypiFCP7UVHnOKrPcSTMXUGYJlU/cU69f1HFwC31HFppR10wj0q7QCED08
DqSvuB94yadKs3ilOEqJ53Q4EqiTC4NLzDsRXJ0W2a77sTov4MwlkcqozUAqPGdh
ytWDAAcLw7TN9GflFTtrLP8yMIyKcAF3N2W1m0R0aSXsczIUT/alxbauM0F8vjvO
2h971zVvvQpIgEEca2Y919JDATecVyJhWSpzlcEIzDtg515wd7yuBKC+00T5tZ6T
aVKdHE1zBx0GoLMWpDiwLmGkKTjiXeEmN+28rSFboy3wp4Q9MmZzSVheDajdvjrS
YVOAjWoAZwFWOoPe7VgBbxzoaiUZnEyKpkSRSiqAqEZLFYX0RnuYqQBjdeqhypdB
q+DDX+D3JxALJu4S8vJMLaCKirfew7I+d5iTHftN6D1Y0uPlwoJEm43KkNUW7Ryc
i2cL+9+p0ciqxi3a+t+I+Jaak2nUueN0O4+MkjdPtkFt9u6u4y/fKtjURGUqSDyU
f5L/Sq+KRn9gZu5LMYW22tKMXOK1Ae8ZvIh6Nufn+7ItbDjAWCzSzlIiRrrYvxxG
w6YClER/lM7qn3IY8gJRNB56K+Cn5SEStLblN9LVdgkjTi3R7lRPd6vrECVe5Hqg
COdOWeW1I3fD5mhTGAY+2o9IWQUtXJ/v0eAFGJN5MEARimB1oyzeADQor6xuHnEV
uHZ9EFETGH3qNMgxR7ndUNIcF6LMst+iDyQY90xWozRNH//7Pa0xtCb8+vzy7EAo
Ya02zeE0iIeg8mDbQWcN0BXUuN7tEc/C6RrivVSDyqCk5oaWhCXMoXt7ueOOErSZ
gPNAIDXglWuTXWsqcktVdGsCF6s5igEO8dXz14qyvvX6n/GAWdejnxGo6MDdwtWC
1izkXOonJ23g9HScbI8HDQvuFFmyPC3hzi2Wmlqcz/UmlJu8yJq2lqXOcf1enavH
42EXt6S2wGKAFPCLbrwvCTyO5IlAqZ2Bcr5iDYTcdIBdrEAV7Dm/LEsPMwavXOTI
fbmk9Vzq0WKHFtOTcrdOwZXeMqP3qa3Hx3GVbqjIjB9+yv4T3bzsFoGLNtZTZYmv
bgbh1iegK9VBaUmFkOFAt4snDwu2QXB+z2J2PSQyQUIBVVMxVm31CVlaCBrZk94p
o+A8hctU1HTlXtmqGwjoGCBwCIZphpr/lf4Ihi2PvBUOgQoBS8K7gzgl4xCg4Y04
zZXnX2/Ls+K3lL8W+2HzSxEIghnrqPLeO36UCJvRUkTs0PHELWI0rimHQoCiHcuO
8kEIx7gjpM3P0tEaXrVF9NUdeLmE6jwCSgGZl4GIuXLujcnjRjcPxc7BxfbL3X0I
ilDmoxiCkCQ2Zw1F8X42bQIgm7+RBjMo6TYu2Ji9anjdz/2ExCQNSZ8Sk8LUUCpG
ZkYte3qi7p+EsubJk+l23+1aO4lencBbrZcvrDm7qV8Wrlsx8VvGIpEQIrmHLYAV
H3gWa8WX1/13FxW44t9D8CCk3xxJSaqnk9hvchODsbnQifvV8r/nDatixrqOezlt
Vtwic84ym5GX6VYuy4KSrPs1+Uv64ju2TgDBdj6nhUTtqtLI+M523BNq4Xbyf4be
RlqtQIa2KN+GofZqY0bvrjDJZeNE6rek1p11mx3wT1t5kBwgyonuozLjWGoXaSZI
rPELM9mlZyo5sOkI7BON7Ma1zglqWqg99GK9njo/ofwsy9Yh6TTJqoz+mT5voMZ3
HBKGArLjBfOK5IT1jWFeQ0UBV7SvGDWMyiD+U2+qAUPfKngKJ5rH6rNZqJRP96pN
QHCY5nN7cTqY9BmRj9p/TloyO8R/t/Sk0lmDI5FXFWG9nHLtqSxVgoG+9AN1Bzc/
RpbJpV43njkKU5mNBeJ5+NeTP2kEJec2LTDUzJbDLtFO90r5QiUko5JlU53R2lqe
YIt7nTYwJAcVstuWk0ASI5CYuD5dUxya7sYqdYxFYspZd8PxL7z5ozf69jrt5SnO
9ZBxE9UuA6kLKsHgBgnFtBOLdjuvuhIhwD2qBPZDBLJcJKwWl/A7cM1r/ybITrjA
U2NccIhgtM1R8LZOJqLmiBjk8lEz/lZhhKTHuyvaCTlFcJjEO8/En9R8E4ItCyAu
gKJTNl34xI4yCf7VUEZijhQkEiUoC2juAcz5Ic5C98qOi9sJmncmsuqB7ZCkoUFU
Ewyopr2dv5Or5sQlmzWS2lIkEdFxspYOb1GPoLXSt0XwCnlDBYy1SjzoGbaH6gLY
weJ0H5IAf9hcfSDqSOK7IksVxwqIy6uzybRxZ4/mob04Oq23KNiVQ+8qVYes9hzH
rMRD9mRf2QrDS6c8M5t4fJVNwvFV3jT/JLaboyECiqBPaGAhBinWTNrxE/6F0F86
4R3lTAPUmIX1xm6nJ33heoefDXqdVP5oW762czZWiELp2J1ih8xOe90xJ3++iLK7
VCPLn6fWce8UKeAObVlhfP/uZaSmss4ICZFDRkPSDWVJyrsrUH7uf7ViAJRdOa+5
Q+K6WneGXVlp0vZPVoJ+XwmcfmZtyaR3OJeEMAZIcDmqvIhG+7WwjfdjDAKSUIjc
PBcWteEHWd0RNjp9nW3npurG6is4Z1cH/lCOnfLssesoT6LV56vjROd+IsGWRCEv
sbP6WQjel/xPJyZvugyPm7kNcjtVMWbt16l2/GgFF/sCMTVrWWzKbwBzz7UiNB/b
LV6OD8xeVUUcaLT97oSGzT4Pn7EKPUmfXlhaetes+gesN4dpInwsbR6jpIDqO6N/
vwbg1eLtD1vMAyLB30os9OtwzzBcoTxngSo21RRREIXVlhOrV0ZYHndGIZab47X0
n6mQJyvIS7ueeDv7eWWbaly7HC3vz6PkQ2nR810BVQHhvO8+qAkFWCzAGuNMA8ng
D5ISZCmonRwn/7b+ZOI4cFLCe1gxN/RmwWW25ySTqWRr96/jUhXZU20wyKspOhil
NYftCSjZT4BioxhpqAS8shBZsZaN6DQJhAJmfXpH2/8MGk0duNUhrDSY7H68xO4X
MaWEHLv/JbJf0q3Q5W07BjeoH6uLu6sbdWlVvFpp5a3kw9GDQxzm1EpAbET+qhUi
vi2FJb/WnRt0bXSs8mrGKxMvbgug3sS30O6rEwbT1u0IeK0u+vQQOcV6pHuV0idy
R1Ztpms1mRfrVNnJ1ogKCpmSKj/cVF6VUayU1fR7IU98hs+tgsKvJqVYouOfChvR
XSWFe87qVM7nOjTkE5xxjzHkXGBI+jnZ5KoWEV4L3PW/R7Xsxrv6rQqb0B/rkPB6
XtYFeDPoKW7jd4GgGzc+CPT3f0ehLcop3mqlbfkvIAaKuehFiYw8KiWsEbQfeDRd
JS5vztmyoGyJmBo0+u5jYiDTWsElgSAC+JRfhmVtZ7Q9/y6xvkSe/7/y8EwuEmHX
XRomhNvm5A/nAXmGnLOwPVFcVjad/TSkxAMZ/Y06ZNhG9yR9XqwNaeseWOlddU1R
tjF8JsdHjB3CD5YzwQQeNwHgjy47+Lcc3zfcoIXXUOILc1MaJ3KoAkTUkV9BNMZF
fxEcKQkcX6ou/svoVjtf40MFMrOajYKZUghSU4pZJObyXNbGlwiglb4xp4JDEtPE
ol3o+yRzeEP3hVX5eyflTSZ7y7A/KV445oapsspGj4fxXrIjOsBPdQXDqitLNdTC
KCKxeblaWX8dznJHlR2IFJj4Y4b0sgnliJt4BtOmwUS7TC+S+RxSTr/ApZ0xu/I/
5Fz184NJi5URfZVV3VxIJi3oenN/LmdBPi3saWOqpIC8njHfjO63PkPGx0Ri6wQ+
9m2qB4UsbtPXQTwQXuygXmMu54RaW9olSsO9wVSyZaDZ5BBQh/KJoxWQkCDKBdai
mi/BAOBwtYg4vAXJ4JsmzQ/tH2vJqUelwdJ9zot8rWPv+l2SKqEB/mfhcsj2JcRV
DU3OU2BI9SN4BA3pus6n4EmsuLuCD6UjrO+dNsZ0BIoUT0qP3aIAd9SPhCyGWmVQ
SvY8IHePZCsrTk+YySlr1Y5Yur3m+Qlv94y6a3X2DWV4YTcalQJF4BhbIJ39/g+7
1Fle4WrjiDlv4+uI4J4eEQBuAGSpBp4Z4f43PSvQzKYDfYgDa/qu28eKKoiH0BEr
tamMol15mw9DCy60/h78gEgXdLYUC3rOx2+Cf689LUXhaCw3LpztUXBErAGsVFIi
fgjt9a7y2MqFzq874gCDT8o0qdVPkuAQPbE4YnDHl9ZZUNutabjfAmcCw8mZjyDP
bYTrd8leiS0m9gI2qMAcqWd5f5PX1TlVud9aIbD7ciBka+AYc4BEfO7Y6ArPpzmv
dy4wlof6pvCa5l2p90QOP4kF3tYGE5ZtD4WcLRYhkG0ECql6aeCGAEicZeAVwugR
Nnr4JhXKfy+lohwM1X8gL6PYslGcqDHCvDrCa+VowEs2IixwnSM50BAzJjUoKkPO
yzaEbePEoSfCwP9HVbd0EtD+M7jbCcOH3g8mAje9Y2apjkqh0UE8QrSM0duprTIK
pBDB7mjuvbhM9VIPyI2CY4Ju7W3475PDDVy0uprGyuYzIo9wqeTMlAoJ5TODP3j8
YauBIZR7g9pZpkURBTaFR/u0eJZWD4OJCwIQ1tGWZWuDONf+CBW1w2ci5VG0/X+V
GY9b5jbaRCe6421lfChKszJhnmLAOA+PXYC9Gc8bTi//Si0EQ5V41hHbR1wN5ffB
nmjTZV5WBzZKB/m4jtuL8vanu45s72lfD211HcqY3sY3IUaeY9SRhr4RzTFy4akZ
k2zwGHsQBmS4AOxtOZ4nJCA/anUZdRR33EtyNn2ZqZk96YkX5EE7J/EMrc4dqTLW
q47ZscgxgsJwv4vE2psO3/Vvrg5wip1x8xyYVsFsZuKwptvJzAU3hn1md7qogXA6
DJl0gG9bRCe/Hya35TZC90CJx3bB1+E3mVsrSP6WxAGddBqTV5OZK/E7cAR3NhVG
hy7gDI0eSMvAE43R7tN14Es7IqKi6u7wxwBjaVVf6vE62SMyNcQuez+4pxOFctxL
Sgi1ZsDHneo8FL666h1F1HMr9z+zBV7viMdgHh5iGmmXk3Kr+QrNU1MBh8wNR4zH
gcNyhw5RzSKvcJon25SQDqRqn0DNF1frKhiYeGLp81aDMmUBdQFFGd8tGfJwYuaY
eptoHWAqOMZ6J/S/cg00beTPZ/qLguUO6ZNGBoN6N8/CXTngqpLZeLnROxDIXH3m
ihbNiJLuPl6jmM0M+c9Nyv9c7VzOf4FhQUJXBSXVmLI7qJlJBoXMRGvUv5+ucSQP
6SX8FAGOFZ94IKEuXqbO+0LPViQGJFnmwCtWosQgARw3ifhxcYiBIjOGON8hznxG
GsdcCCaoGgkpT0WA+DTU0o/nWXI20QMHRyuB0BFsd59M/ego4GDTvI5AnFoGXL7r
qf6y+J1195LlyWksDoasVQAgru0CZ1ynU1S2PvM0OPk+m2asH0YpeuUMtYi5h2Hm
foVPV7ZhRK5npr+d/xfMFqZRCGDAguvV75tdI5P1Os7PmXpQ7ZCwTRariqyyqMrW
lDMKag8qfIRRIn5C+zLdokLDIPxuiTNK/kmU2j51PugoCnUkcs1xjdAjDGJsp83q
mL6MN9fhIyyCT8nD2bKBD9fLOVWOlUmzWbZRYGdmJaQwUUE6Ue7INjMu7RpUemhF
AK1unjEW3CvbDArTW41Tma5jDPTg/00fSnZNDm/8YzpntIIIN9STXe08LgBgZwFN
LhW38Mw2Xgo05e2/FyYpjR0PCn2eIh+Xs+SRR1Oohz94UBf1SjbFLoa2ssSeFy0j
TcQj4WJPv22c164vQD/1fSdbDY6tQ8saJrM1CnWjcAeuQymq137wxhRXmMAXbB4T
8GbEd9nYwphLml+L45RSIEPhJn5eqgt1+ei5XGEnL4tDtigpZeeMTCaVNRPI/KpI
/UHZTHmGgHP955KPoEzIv5/0s1SOsmd5hNRTBdDTYS6z3W2X2JIhKBH6e9HYx3Nc
vVXn1FN4q0vpG7vuEcmvWcGKzIJdzxOnyFVieJAKsuochFe8s6jyn84mzO8cN1to
frxh/L5+AqrUNmeK0RQTkvAQwGo1oKGRnl8t45YL7XOgZi54kfEpAaNLoE2cAmK5
3nw7Mbj00LY4Pj2P88aX6MrQ8gYfgSuxvEnW2MqVCbXC3iLOZ6PEItyQNHgEJZBa
e7xX0iigZdP7fGoMWvVrsX4l81jXzkjtXBWJvCJ+6xklhRTuX7BhI9HAlsLSnvqa
/uguJpIIJqyu1+YNLG0CuafmgW3mToLgxRL5iyZayFtXkV4sizUXjEtMq6PN1gGP
gWuxMLtEopDIBOE9Vc4mP++oeAFDHPHHMQ9UG/t/WSTHdPyBSbPWdNvnDlYPmrzS
RdWTgFYNzyw+Yo5yAgnchWOnMWltQH/+gLfsHavZgj1eAnRk02NOhkF8h5DPvBQj
s6l7ysZSDoz3wBsE/BHaQiZqXOY5OfywwFRKZ2kjdBVBN2gLhk4kJZ0QP0u/P+kn
Y44JSOAOJFCx0nNPtoDhSgoYRUmeKPnSltr8I37we7qzNVEL2Ct6ZFbmWnuU/Hwz
YICHTHj7WRlXlk6MDS6T08wlDFE5JV8vTP/EZAmmrzT5sc0GFteirG2tJk0mHtM5
uNEBi9ZXIp6TxMA0TTSZiv0fM6tRyz2iksAz+Mw4ewsV4+E6hJMVF8toLShofXSR
wTqU/jX4rZy+Nw+7VdrQDdHx94ANBr7iMHVFxYqPiXsmenssH3O96f7AVq/XCIuk
AGMS96HSqEx/KT7NHO+Dcb1LoawhviDmQgvzBJnYhxTd8KauqnsoXfQUG9R525ds
R8T8mksNMN6MQlQ7T/xrG+F5WEi9Zy+E8r1UEDUI0+ZBSp2ahCcnN8WZ2BMZJpVa
7NapX9RwRPLBNUzR4XX0t6I2YbliAtrQKLcscFDJObGNyuxksRnad7+Hc/mZdVG4
fyfMgSSqeHwzs4vl9jSf368zgBTKdv/FtInPXbf7F3qrEMrn5MevOWNDbAp6r/fE
F/0/XvsoFUh3WJJzaPFPjGFkOpIlRu21uNiR5mxCZlBvNo4q0Bzz3X5bFV/vrBKY
QYyl7jKSmmxKM4XGXHHt7j2xY/+z3ubXODMaHWOPee1gY+VulAj2U8Lk6lbaGeUd
F3RihQmINBj7V+9npIXlXrw2mP3r8ppmArUCRVD0gTAos+pbS23R6ZZg3kVuWxne
9XfolrbczhzU5HEiZ+G4rCSMVK2N7g98ZJfQfEY3vgfmryAnOn9bU97is6bA+A80
qnv3CHIUYtIQcB1Qy8aGCYPP231QMTETZFxTWib+JIIMy6elVMszIYry+FF0Fcqq
qu42dOtBvKaDjheoE7hhQLX5X9nljTp3ULlwJJbMrCLjP6qlHIN5mnve8M/rw8s5
MMafrtE6wAURAHCQkn3HyvUd1OD3NhDdLpN3xpvcBfwrZXtRKJFb+mrK1R+lLXQn
b6yDrldXr+T1a739ykbOx554KMufyfVLOmbVS2AQrv5zineS/FVRGkWI/DHSQ57E
QmSJvxeVKQdDPCkjZZ54X6vzxqCZc5dg9wiRmnyBcVJ+rWK6F24nmc2HwcYYcLz/
odSFRkAtirK7gAIS7KT3U9/H8237ATFmNXKLC+Q917mlamceTtRpHdJ2dnORq/E/
HOu3pZdzKaVSN1szycXxAEXK5OLX9LuSJB0R+VFSYLkD83DgxTwIOpR4sVxx1gVT
QlWa/AHw1gLTcst6QAQ/B98qaf/ZZl/yrj6vS5szR1bRzzFq/QyqHfThjMAT1Zm9
tcylf9c6zYEDbjedtIOqpyel2noxs1l3FxYXoYAQU7zLU71GQ/HKMmydow6QIzhb
zDFc14jLwhw9XjT3BIGSZ8FsMp2NoPL51gympuyFqh3kdXfxEJ+OvoGtN7ud5ATo
0joGT+XMwKKgOGd+ZGQ4hSU1+l5JN/G16qAmV8tXD1vpdDhY1iU/8Zan3EJBK4vR
rM5t4hjc5DPmu6NkAlmI+V7BwWTGWtwYr4X3qRpsmx4ZXzrN/bvyQaOdXA2efmMU
paDMoQuL+bfQYlQ6ayjRWdn++N3D9bhGWeYpnX4vQOnH5OzpE3n8ebDZpYf65yHb
OcQbGoDFHth9i98pgCmRe19Zoeie6puNsmhFfzcx4S6zgH5aSFLJjkKZgtE6+V0U
a4zKH19O8YDviwSiefSjNUzYJNOy4wM1NvBAjVbQrvD5rJIrDF/I9ux4AQCr9zUH
0HdEXWhXDUa25jy1hJ9SF9nEh2pjppuaAXNSABp1C9OnLA8gepCuXXYPFoVqipYT
xYMIjvLTWwrISpm4jcPw45ryddXH0mpyWYpLlY0pNGDaWlin2FEhYlr67G0XOPu6
fbLlDb5hGIlWSq155LXI7OSkcjv3NPbiT4BeXDnGZtG4pxI/ehYF4JQnO6xzXLnn
VsbZrsQjublvM1o/047x9ispNFphlLeqqpmKcfTA9xdPA6tSVufiXx9F3Q6JBy3h
mFfNNe6qgZQnymjb+Lm4XGeY9IA9j2opOiJ9gAaAkp37ak3EkftmDh+PyvgzvZtL
rmuH8WQgRe5yu0H6FXKT7wTTr6ZbFzH2ZR62d2RJpTuQBAT9zfmXuzJR1gvZC3pO
wR8/xpinrHu1pKtKiGpKEmX/iMw/cYnkHgRlUyLtFWogqWa2XHCpb94nOX5Vrjy6
c5N996NXVHPUPUBPkwkQ2F+t5XZlOytoS+6gdc+vz+GUMAmbT9ByL4XOyM4IR/DO
r37sUJ+NWu01PdCxmsZ3BpuwvkOaX9Fy/mlXu9wOqk+A15V1zFGT/N9p5QWqAG3U
kiCH4z9shxiNAqI04jP4dU4EDqzMt0hgdnkpJWlqVTroAQ5N6P4bHn4etAJMQsYT
ohMk4Y4rq1RwuG9nnfFSNLJf5E1ArSFV42Kx7VbzzvdJ9v2hGNOHKfK8WAbX/8jb
djr5Oly/hR90xaMgnxsIwaw8Ah4CnK+oaDVuyU3d3o7U8mYW6xx3InDe37hyBfNN
xiy+QePiTOixryQ0lWobxr4aOqr/RyYwrHy7x08vklckLGxSRqLlgXyRm3y4aol0
yOp7/B7PYsxbFvahz1uokgUqs8uPSB6T3+vuHkbOpQhcCarnXs2KOqhmHtHwOC6B
1pM9VGblywqpJwmDmnMHICbTdllF3bWwsJ6+3B1UxerqIQ0/BBX8B0e4k3ruMWfa
BwIIPoGg8j6pGKHRT3loYJu72AQET8pKddMo9a6BXIqH5BUZshIzuAbx5RkXJ2Ks
3P8LsbL1fv32f7qinCGtItKrYTfx96jkMEGsXDzfaJXc8ApKYy6xPrIrsCYUQ93/
BI+cUg4x6RemGH/w8f7ALZj8wRqVZZOazMLHVT4k/XOztOR8FVeq87+4KPnKIzwh
RLnJMfTPhYFFU6W5aCMFJBT7j9nRd35iHYS1Ue383iTc3U0R6aLQ9hrtQVDrT9T+
xgErAwftipcCnVcDnwZZO1tozNYCOJLizIIKKXePMwyiVXifBTqSwPuM9FuqIgJj
dVDRpFzkngQdnhOHtezpoP4+EKyv9lDO8vIHSJlOLRa9V8FKiY4zg4wESzJ4jJq+
UHUhLt1CrSprzPRlfIgVEvmzJrOztBEyR6S/qG40XQbUNKBL1sMSme7F7lbAYRn8
GIo8bnmmW6fppKX2f+Wj21QQ+cZB9Ud7e+ehthtGUkJcVuBK/keXlceiBhNvEKiC
/3JGIbkNXyVIPwuqpvTpgzx6ZVxq9nIZGKLEsFLD7axFY6o9biRO2fl+fAvVW/3r
GAoIAqMIys1q1cTyDeLUzYlKeqRyCdLOytdpx5m0vvUPbhWyLk/FK4tNsARsyMRc
rrMqayCWcqFHR94s4rV6CqzAZxkyublucT6X8uusRS/RfbqFVGHTSjLlePBM5Otj
WlOVa1Ito1+Hq9mVVdiL+enhcKT96BEwWaD0hDoDhijtFmAZfT5/pysSi1W3arSx
Plna3WV/ozry+ZpQ8t88n3MK00NxeD24T+o2GYBGW/Aw9q8N3wi0zFv8Iy6curQh
GA0pAiFQP53jCnHtO4J0nT/QATKPfhOJptSMRClv99UXR1pmYMkSCiH3Frz0cD0/
3zb5DMXIJW2PgJII0G2vPv61+U23H1Q3QdcJHWs6Dm13YDpB2+ifuIvSgu5mGNDy
0pPlg6+I6k7DNcz2SAVzs6CxIAZc099LyaVBMAyHGhrfzrr4D0BMZpYmKsDiovN3
IT4WKCf6RkKS/X3ybjBPuL7a3VIKgybEnwTS9Onofljg5hxo/iUFo2gcZGT030QB
32WmcJyfhwNucYu53JuYi2Coe5wfGjFy72y7Um0yfuFLzrt+Am6vs8Kt/D5IypSn
qLKLkyXrREfa7sMjPg4NQKykwTo4a47refAh/iFAhmSSi2XgQLk1ad9HkRfWyIDq
tO3v0eBct/Df08Gu7jRaPFoonnoajHrQ36z8eUyqAzX3TNydSpicyWlQbTUniDCW
4JRPmCZuosXrvIqPdXMIlF9vtPjggtbZQ5yEDaNd0TUGidCtGbaRgoocTaIRAAMz
eU/XpHrHPE3apqNraA/axlJ47YebLqNREbHHKEFHLPAgDJmaBxg0vTfHe84rghPp
/wEq3ef0nEosbU/QxSoYS6OhXm0Pi+4C+jQ/iqYhV0d4L8ua8afN4xmuE9uWH6Jj
qH6xbYzYcTcd9Fnsw0shUfyUUd/dq6tz32UbOlsBVRjZFvh3IgI2YW/tR8qBKonM
aCzzqCzWyzEJCbTnVzPYYiRhh0j9gJfKx84DgUUp9cF1nH3dt82NsbfcC2wVUv/+
OAsPqzCqmgl4X+XIu3Q9aeXnuyCcVAi7CNKjrA1alYsPzibxzl684KG1SB5cLfyI
Yc4OEl5HlHchEl2uN1FjqnEvXRdVNRny6Z6fbQvMcxm4gKI3zdI6c7oKpo2ZhXxs
8YuydNcyRQoIFUd4fSoLFzcliT0Z3UXBAmJ3NB5SnbU0M+KWgDivi/oArQ1aIOYF
WAq7fIqq61FlZJKgcwb4QD8haMz+PrWqHeF9PwjzH1Vb257T+5JS3yk4ZNdMkdSS
ZMj/hkG9i/P0MkJc6s7JI0OV4tXLENnC3b4uzZB4YlfKVpKP2d6ymRa680K87BsP
64gjzfagMN8+0/fBl42sMe6IrLBO7OjUh3q2mE7oBUJ1uwW00sy9u9Q8m1SJUPdk
CI/Ks6gNxZlxtw4kqrizrAqY7WJmUOa74CyJM6mYe04l26oNyENLvlKo3MIptfHN
Gc//zC5MRuyZgt/Zo56pmaIuv2VVUSjjjLMVsVjP3FRArEPANoX+LuF+/PF4snCm
3Nei5RiHqueZmxpKTkUd6A6ZWC3WuJlQxr2PHAlDuHQSZfDTaFh149visBMQFEjC
G1ZirKTXFFt/bkpZNxmMsFgrhbYwrCJ42eylStIXIr0KBJlzfv8yb4TKsOSBj9PN
2qWQSMMTDDIAj91AoO7VPUTYoNKC+nwKbEddhtnCjBUEyme+bIBSHHjlW3avcnSm
KouqWaTW+dWwOVAUc5QnjHdGGe/P6Db14CnbUf3QvcjCnNiKooNds6FY+KkNZY7o
OsYHv3Ydu5wSQJcCW4YOahkN5pbUnP17yhoQeuGVtHULBc73WYmTyO3gylOo3LMB
0NNqsxt4Qn0Lz2drpMtOrl4RqAE+aeaE9ycr+kFxFuajBC/oLA0qoV92aNefI47K
nL4gTrOd1uEAlC2XndbqLylOFOINrW3A+Fwele5euDpL2lUPdOIHe1XnOLGfRUSS
bTLtn2D2Xih5ROdn5HvYcubyhV3qetOgWKKvf/FcW8PYwabEgLsrKkvMnxpRg731
eZiKZIhYXts3lhHcT8MDiamxvJ/F+SOhqOpDMQipmrJjIsEyCEz5ODASZ7HIH2hf
6mdKz0v7j8rNb4WUFtpC7l224j6uiUXG8ohRfXdhfXwPJM7M0Vz3VAYeoVidir1m
EAGLaysoqvjZrMy40lOtzVxXmd5p4BrH6y4gQeVDx8mp9wK4VsHKnjSHu47JMoZR
n8Grhzw5yXWhTlERYmwXOFsEoYsqq4PRuj3RR1ZVzAB3ngWYXvgTu/F+4h6ROGW4
0eU58skKSFGGyvxAw8kSJH1gwXwttesOhB3Fun13trXn97sP4X+0pjeX9v1kGUfz
I/GMMODSvf1YZlpatazBxz+sYTFFvgAE1S17Vj3Pbuvbu/bKhfwEmBbjlQRvQeCJ
KUCCMyQisX3OrJV9kEfHw6qOibErL/29gRW5DkaBAIlgt/1SPDiGeClmSGOqFZn8
fMpmKo3covzkeUkK1WvBaEyWgpqmwRmzXDlWC7XCCFAbXTibbsyj6rpNaJfLXEEE
B6K7zTKx2JjuS6BZeKYVOZhe7OyV6UD+h18t1AtKrb3HfyGI4WVWW30tx1NzRHTz
PIwFqeqsEOw85+rHaBUrmzzZ5BRqjDUPtMrt4QVIprS95oQPpBP+UiQAOdS1dl8Y
qXXbHiq6YYIAwAd9J3HVsJoOX79t2eL800sgeon399qC6jvf1J94G1JCdLb6mPZq
LXCt3e2+ScnuIUafJC3feO4mjRW1yx2pE6HSCKzIFJbn2Vde6++88d61iccX9CSr
wqfmAegSxmEdnR08TDt3TVCXh16U/OOhJguR4kYDWlK51rBhBIK3ANZzRhUr9KnY
IrwG1w1UUAR5uiO4LKez03ikDWCRwJ/1ko40OuxEa9rQKyiqEO4YcVyn5fnFWiT0
ft8yITt4vRWaymujvcjrtiTh11SAwWbn9O3yFHCLFTP/bN3XuRL+crgC/UKtiR+k
JF/phjuhlKykYSQLzEzzVbiJjxY3S3MN5vS/Nlz++5scRNYrbzCE01HI22W2eia8
zgJ+muuKmU/Ctco2DwZmx7iSwcMLb1i0WYjPXGZ4ixHA/AeBWqp6M1q28bjPOh1c
OfnswTAb0i6uZrrGKXxmoFb4tBfxc9mCIE8I7l5nNwagWd4ssTRq6wgRYR7IaUJK
5vFX0gP5GiN52qv7Tm50xJ1CyjqsT4xwltFrjRHDeLE1wXWa0acJ2S4NQzbKp58c
vIwIFGecQIEaLcAKgr7O6emLUtZhWHpf9KFGk3deerV7NPr1HPc6XagbBQee6x9i
a6dRDf7OAuBRJkJ15F7IVQF3ZrShe/kwGPk44qIL1lze8GvswBQbccKoiQArKdQb
0qYU123TicVBQf128dSok3hHbwCoGjPexyuf1gK/Z80m4gak50i72S9/ccZ7Cg2F
KxQjFjr/7DwUeezylU/8XMQPbfExnuYYc5UAr2Su+MOjG0JyUsTJfCokztCXwshi
Crzu8qk/EqJDid9NC+Aohw5xP/MyAjWrDXwXuW9kHbfGusWCtYriY2eOjvtUCNhI
/2Iwk5QLw/vcgLGGYr3YsvjVUydxrdlKQ29wOJhItO3h7cs+6Um3EwyGciAwOkDw
z6vMjbc2i6bhCql0+A+GbE2dn2SLXIF45DQRsuq0uGaEZxrC1LenwnD+3qGsUt7O
p4cvcykVpnhnFqdg1/fc4of5KcqADzb4q/Phd7tM3RLQcKLOAEOhtJZkQge0Au2J
J7blYQ8mi3tkuUk/6AYSjVracZWhG7z+vvfFPIGqYaXHqaoA0PCLvNCCQAMp9QtC
2J7I5afba20wDNizesn6WTruEL2f6kmBefDISXryGfdT1RWyo5P966zYC/3pM8VL
B3SWr4RuNTTCa+f5OL6W8MQ6SRT4VskENFOv5NDTpPLxBNLCj1U6e5vAFmOcjE+x
uNSJQhXTArNt7jHr7yMly/tLi48PVJs8+OORQyN2m9FbnDXMBXZEYtwS4gk1OFyS
JFymRhwOZgaGlxC8Uhh8vC+WAYrIrzf5mBfYoipmCh/r7+p1Ic0fK0KUGdEGqojh
sz5H3T+sYN59aJhsK/lpIdMZHIQm8enV3ci2QLbjX95UbgFRrQPGxQ+M6BiVQTst
O2JTjlJ7xxqta98EDFrK3PY9yxfQ/IiRvo8gVuenM30EuuC8lJ4v2rM733gOwoE3
FCTCUUiz7MgI6+rsv2/DHovRP51mlM5usdyFCtPeIDcBDSwsJ8t8Jwsjjp+RFk75
ZfCw/zI+cmnVwqo5ZIO4Ym26dkWs4VoNV4YQuHpXt7Ola5mHN8qr7e0npHczAIK6
OkdAzhrhoSEFQ6eD7W9rAgy6h0Q9TJ1C87BRFrd1VtbQc69hXpnQzOWgRWJoepaO
SF7+ob/8L0nxfX20gav9guezROwtyyGKhlckRGBQm3gK6IpElxRiYePBfPOY4n9/
FeW20RiUeAKYsX8BKiHi18W1vzeJsg13ctYAPgjnXe693dgTahfbjNsopfheVxPc
XZkiDYbw8SAbV+hrinRqhsQ538Cqk4T+F+N9895VFORApsxMxk0b6tIH8pC601lz
ExpSNQEj0L8O0jjovyLVIYH2MhtHj2Iy3dQWQcKYkqdJIC8P9Pv6PCfX62CPH4cs
W4cUgeKuzeLL9xHEUYs3QdzDYjhr+ijcpDwpMMrfTEcpdMoRb/wjkFDw87UNWcZT
Vc/wwYQq1hdvGoUdLQ411ocNV0MngxLI4eJDfZPLjleLaA0tEeNhNWPD48kzkSfi
3xqK0zFVjTl0rOVvxe4fL2QBNlw8+Ms1zw2FTZiV6jzw0NM1wXDWBTn188hRjj9y
ZPD9e0oGfeTPeuaJk7S90Ph4115kQxrZDKZ0tN5NcUtJbRZufah0wzYuxQxhTA6V
aevcPdowb3EdMpjF2BXKV6RX7qwNtvN8aH1fnegdGWvAf4ldEpm5Thnyc5SG1eE8
s93FYgrBmsWRJILkIo3F+mUZepUaZ1Nkqag8PWhqCZuo0Z6wPH8+/bSKn5P3PrGY
eL0hBKBEH1mQyvXsGIAXTcAWeZnAv9aFChQ2VgbJFw5WsJXcNbLW/kCYLE/rSK4V
Am3mql31roGTumsv4OhLcnLuGjjlDpKsWmGjRHO7Bzbbk3HLCfuDQgf1HZnQu19o
9rJy131asDrRvRVCXpoj4uYa2K3TomfscFeeHZhPapbwGuPDqy6VfcJMgF7uyjPY
ENiyAzC9C0n+q9wjzO23rsJGkUj63VjR/QyKQRvpEzX4IiBJlJozfzR3rVqQY2vc
V8esReQLwtIBKjpGE0LQbu4XwkCaeV5Qe0zGkGk6YsE/14ElU6f2uRIBs+9+kwty
cU+5fj4l88h3MOn058b5cIC6fLI5iclLOhl32B8OoawMN6FuURhfqAO4cbXXYsvg
6CWWz+SJgrFv86W4oQWRLaSgDkuWCyRyXnZamvRPLxucpvJE9AYoLxfg2j4xpBTj
ewtw4tdhiFXzNFSWleDGnHKLDqqpa1BoRMRzcZEBvFBuNYXqVtBoOs3ms1jD7xRV
4ny3MDDu5XUNNMtIGooBe24jTuRbdQ5t6/XfMEJ89r68RNWffD0OLkwPrrpGtTQz
lxIHZ4aYr8SQvPAkF9hPsA7hQTFjrntztIO+DvkSEPhEfBVWz1lWYaqjvndveajZ
7bbm/I2voSsDrdtI3qI/ghtmgDTEwsboQDSuA3bEyTqjk3CPAEoQn6JZe8ANdJVh
k7dzUOEwK1U3m86XOl5vt6gJR7fJANgcmn0s480Mmq3oP3oo8sTk9ZOXVdYhMGTF
iBO3rO+jZ7G9X9c2RBu9Y9NqeoXf+Bxqjza0lf88ioeAwo/+y3B20vcI4pEApTGp
oJXr+ZmyHydK2Jw0PCIdCAAgAyoV/2d2Uxq3Ml3Db+aP/2MhkMvM/bvtBl6OhUhq
rPi6CI8hyxpLo8XrEbCU799A6AYCLzhSUHBOS2exaKCHyxAygfrSNN4x1KT/x+yr
ZXWrJByQJay6j8tO8hUWrUGc9BlBArBjtSA2ZRKEyupXeUbriN34KRBS3TY+P64Q
+nbyg12QPSK5ikMHSizmdbauaZnzAtnAPKYjUSsfI0Toshn4HXWiXM09DiZJQtsF
iIC1kpF/G4aFJ017LaaXwQ2/rt/GXWxqsEiLSkhbHOZuV29+ZwfD52PcS+jICfji
O1UhW2o1FMzYOkiPE2cQatqgTSlAft5/J1hztPyCFIvOkiTWeyFLIh8ilHuDr2Wf
CWvpGTkKCmErgBZM3IRWdu6H5hbBqSaeYkY2iwu7yaGYb9vAXjfD4iI+OE3jlLpP
G19G8GkzG0lugTgn1Ynnz0iKKoMqOnH5ZFksh1lJ6aSCMqGjGlZuVFzwU4h2vdCq
UsiR5HatwsI8AvAW/2x483yftXDlxC+qH0BCQCHi7rZYxeFwsQutQcELJnJPwpWM
DC8VCppFmAH25qt8brV39CSYKuMPndpuWGUYzv9EL1wwMaK/I/TWlXGwZBywkLYT
pAvdkWSlYz9TeGp/lkVTHnlVlKL/w2O9/jyBJJsvMTMfk4B6L03nPZ1ONo8QdhJG
R6ZuoeDyqiAdGVIic1OZdJ1wrvo/ouUeWlWEfPQngDyoa1n3VwNP0LWxLCJCHVDK
m9FgzBWy5a79vUyEEqGqskLJTz42qbXpe25OyGagjm/Av7I1ZxUYPMJ5R1MQoSFU
a0rSWhwwrXjNAu+mMvp1L047ewg2CDxJldLuFHl281j8eh1qMeUuhbIAKjtF/BdV
/89qL52hBaDBI4vi/Y/Uzp0tfxVTN6L71aqEzQS06EKT/+3QK1tTiJIwbggTjDf1
/njiD6x6BO/NV/zZ5FuKGfSgMh2Xjvs+MbdsICXccShcYwHfB3fsvocfxQ2Wh8FA
fbRKmy23ZIHDOoY/wdsJTbgXqvyge9oATFkg4SUF63/V/ysHAvrnBIIDS/l2u7ir
oxaL6o5Y8TjWU5g4oI6YhDDd/O1WKStHYIR3hSehjrBAYxTtKVeKBDWTkNldh7Md
I0UAP+PcZIoCFT3biLy35ZLW+TbQYeUsZQVMGKfGzn/y1MOQi6BM8Pd/Fe4/WMbJ
EHHWyjtFpBRVSFVmUpN4cGZQeD45WwjivmiJ+z2KBWi8P1QfpjEh6paMG+qBCslQ
TnI41UaKV/Yp/tpr20DbIOIE2vv0zUcHPUSx6mvnQjRZiIkT5jLgVOGfIZ4ris2A
4PdzrNh/S1bOATQ08A6zXYxLrrQKAfp6tP3V6uENiWFvDO9j3ESnymVK6P8h1qsM
zkZIEBogGAKv6X8TE+5R0eLPb4WXj2pV0GrFVQ6WZfFvIAUtoAMhl9R/oFGaBtLV
Z7MA92bvl1GmEyCab7lAWxBszSvhDwUU2NC4LB26JlhnsPe8JkTuC467qWu98XB4
N4wOz+kgVgf96SNfrKE+WFuDJmAnYQ+LcNHdpwKKmjvCNUy7bw5H7TsjRIfc4Ay1
T1GvbA81Xwox0qpCRfq4LxyIwfz9EaihKe2zCYbYmlPd1ILJAdvpIx1mzFlKwFAh
7xuzrJOzwasHjbAyzYrgl/ZmobxpIx4LTjvz6MT98HkiRmZGNwVeSvlhg6ZGoNQa
z/ls0UtIMRuuRSBexoJ8WjAY4Dq6VtW/X+YFm3kkVGVtUHOAwKyiZ6OJOCB8aLhm
lUKR77FIExNQtVBRtSeRY9XnTKdNUkwjknX+/ufrBs16kcojf1cdAxI/ECSgDCyX
PFQ2DX7CptPM7LwvCRGas5mo9Y8bb2uENEkMTdDt/8XL+Ga2LlK87znypa2XzkPw
nLqInL8zVz1Ewmlpdc0htPcb1IQ0+kBkss4yDLz0rNdwX5ezIgjhVXqbxwTz7IbR
wIojnhKr1uy4cWNCoj+gMQ9cDCjV0B4maizWQuW1a1JZL/1qhauGBj2/odaHckRT
ipAzbb/JBU0MwMhLPiMRMxmyCKR/LftKJA6C/ihj9Tgt1AVSnWfz63knYLMU0YVJ
aLvxszxLwG606Q20Pl4rYj0RCoZDHnnFiw0+dGtHeh0d8UkLNEDc+5VfBlAWFKG+
be8+6LQRHNdT6q8OdehYquCcP6S7jbObnUk+HW/Fki68hWX5dOz1WhQn3Op3oiqe
qNI/tMVHfFq/wdIe54WDlxqN4PDPxPPa4uKbaqrAst8d5adx947p+yvgqW5nmURK
SoCUD6lpFD74DNqQOtWzWhQYBv8VnTdhStUaP9AL1ctfH6bnHzBdhi4WUyAr1jE5
5dYmroSpf/ti7cmp8vaSo5yhkLe1Rpg5EOIRtw98bssFNBZKT0LYgjgzTcCXpSN/
+QHbcO+d2yTAUPNL36RYTwxlmL+NnfLhC4ILhmjmLYj4qwattVpopab5iYTdodFL
p9keaQUP0hfgq8G8usYt5Ic+K7BUI5YXUENkoYdHxLpGAA26b09wUjT6vj9tfZOi
Z+XMTa7az7pLLz8H4E+Ae8Fn/g68dEt45GxhOrOZNbXiOZhbdTztSMV6dsuMHXCx
sncvyQSwpHNuaH3Ht7Jun6gW58zb/O7tMZzRX6QfYfrDC4gDRetQuPaB1gqA+ReU
fGR/5uLJYIq5PIHzBtwJ1R+kzjmSwG/nJwerMN08vzX01TkvFtB2ArgHfDxpTs7+
Y9UvJ0U5rGitBN2CKUtF7ONFL8ckwalTL4cCZQgUnk0UQ7fZ5zAA6ZIzC+d8EVw9
9j2uL697fM9cJsfnMx9PgkVqa7Rhj9aUbE8hgh4BqE4LiyLgO3InUKcMzOBSCdPD
PJMWVQS63VBfYn5bXlql34YJxb55amWuSjgNkYjJdek0gxgZ9O6nEbD9ooh/AFUg
xX+5NpX9RoecKj8efG8zcCk9gTz/Vorcy28ORE51BaYlKhuNbWZpzURK1FDPR0JN
ci2/O2wFHPPsEmfHmuCYTgKDnLZQcP3rHCJVkVwDIorBMoWzF+Z8PJlIdhsrrIHY
QZNipMSaKONk0RrrB6hyF48pmt1GkTawMK1UOjW6fnREuhoWWvXeauNT34SErIiL
dDdl3oEImsatg+dAx4IFFtmcZHD/dNFw3BVrHEwF3ar0UH7Tg6iTKS8QBMxnvKJU
mthhZMU8ICr1J0xB8oUZdnGfkOPzD/byR2YXOngqtVDkOQaeTtrDdGukiDjr4BLo
AOVpKukR44tnqI6Mi3cYmYW8zeK4tXdY0EQsTUy8nYsSthbNLGo66Olah7P6Lx8f
q2khHNOmUZSfDM9fPrwfE4Er86hSo45fDi2Fv0pVsRi6ga+FS1YZ+acU2i6/F70U
W3sFZjW92GwOICGTF9dd/SPZplCLMjyBmDowpO1rkop1qi0voTbge8Fp5GGZetPE
gPeI/3+0t1+bO3Zb/rbwZXrVsuQ4+vMDNDD5S/iZGO/2G4jdR7JvrNObENutHtgF
LezJo0L9KY3V5m2dKb+WP1XssPgFrD5n1EhOvtKS2Jv/q2tiY0mwdDomcQwY9sa5
ZOiLxXk9WmW2KV5KkwNxQHRbVCjhnpXJwlMmn9dj3qF7egwv3RAuM7HqP/HqfhNa
DzCenNirSDTihm1MUKH4ahiYx6Uy0CfcsXJOo06gbBH/8/nLQP2paKekRrfotjsn
n517Fqo8oJv/9CLapKgff16vIcPebbhtx3l6Pvf6b+pE4yv7BIuxdUEYHsSGzs/B
4bE9f5xhuyV3Ajo87Skr1anFHv8C0AFLX8TFrbRKvD2t2qgzebTOWeBeh3MS8+60
IlyUKHACR5P7OPUsfsCARYPIG03pLtazQSaPPXi7Vv5iUsdM0StjklbEzn4aaG0U
Jl9X74D3ZTY+L67DqbbTfHNm2gigv+TnaWul+vLmpMpeJ9s0ZS/xjYp2NiLzCKi5
JzU0fmmni7jYGpDGEScHR7gQQ4TicvOdtfJH30T1pSBfDWeLPzjDeYXsDXkw8AIF
U1/9ZCg9PXufHsgND0X0AU+c0wq0tCISazp2wG8KLVy8DsZSdUsL4omKXFW5YVGt
PREhnlnlM6tRL1GgwZI4LCg4hl5DOyUtLGHV67yykJXM36b8DIt+2AHp5SACULEo
ZvpUuy/z4aVF61k7zNdtDYY4AATm/4nDIcrVASQJxfYtSOaxwt2y7i9mlwaB6yDp
yP5NvOMMJxuLKHgYgg5hBDC6kSGr6J+mT0GWGU0QDw/UGWGpyeUBeurisAGcctGC
66F+1nVuxEoORGcLBBgVxO3dmQ4q9I18cZm3MzAzs+qHU2VvFW3tjJoH4w4cxByG
MpSEwo9ufjO4aBfMzP/w1tBii9qyScqSStzihKNnblZbno2wP1CyE+4NiarBxf3w
vGZK17wh6dE8pdXIXykYVEgbYuhXrbe+KsuBvu1ueLSFZRwhVUV9CXLvngH9T0XC
lW1KyzDBtiE3xmqic/VrHG8FT3BH58XyVjSxQD5mINRoJZwMVGAPxbVv7KPyw2jn
zYjuUxfHecELT94y1CqnV3H0mnfXBvuaTNIX2x5wnD9pXd58ZyGABULxWPu1pRu5
cbK0cN2g0gvXR3JHLArTvDvJUBpT140L3bubJhBqXU+Mal2GABgKNAPJ03PxYT35
FlraeYHP7eGvdlCVEUnovmbE79HTyFfq0bz+3abxhbiRIZikxKKAwqt08jec19zo
AHyp838Id/An2vvi0F8Vtv3ML7K5ynNPLtPAXwblCsnMeFfRQALAL6zRqroStHqw
qAIR5esD9vDqkfJw3gFeJdG1pTnP1G5xQQx3AADOpq7lyCnVWjzlNq/4hfkKPCH+
b2E7+rDufc5ajTEdnu1FXv9kPn8/J4gPTPugBzssPp2RIcQrlQcaajbVK/efjvbW
/8p9AH9tbTVRyJemxZVn7UZznyU/foG4uTrc24PFxf9j97QGaJuKCzsQkpiLNy81
GME4/4DQpO5Dk6gDO+E9CnqxdI5xtQ4moZ4AJBsgfAuAfS7f765pPZfDlN2Cd/38
aVF4XoDt6NMOSzL3LDNOdUOxcmiZmkb4XckFWaHdIFv171LVEJWDOWlSXSRe1d2y
D7o5PovjyvLdFTwzAexacqXUPxrs0pV6Wup0sgo3d1z5MujkyrndI9GF1ptX44bk
Xdnno8l42UhnaDQyaL57YrVRlY2+zPw+gWqwoRvgpmOa+MORaVh2tSI1VqhQHXWp
2/SR5r32ZdegUOvtdBRLFS+V9AdQhG9iHL8yYOSfByZOqMFRgMfEH2/Fvxsk8pC3
eLPovOTjBNQOcu8RIWqv4ePQrtPhYh+E6+ZpiAqtgQ07RRAP6cYwlCXnum4OrwFv
4/hHAXzWh556K3u0CkYkrgrPBNr3LGQ0yBjnK+fLPKs5yvJTG7QJLYen04XrL+ee
hmmY+eMilhA0Dg9yOMYVuFX1fK6iw2qa4+Kz/Ozr5KtzNpXIUd7BqCGNa8N68Pao
pkXetpmqdseyEm8Io11b7NpVc4ql+gNqUaXsWro/2nP9SgJeUxXU3CtfCjNyoK4S
GJXTtltaVDLMJqEgQVqiyLSsHXVpfFBndyb4vdeyVrSFFmRHsvwnXs8zHKQZ78pp
0AcsS0duaEZzkOIdwRY3OG10unvYpaDdxBGJuaK2qNklm5xIuUlYcUwhPKoj7m36
t2JmVXpi7fcmJxDgRmye5AyoyWmRm5YMRJIc+dBH/HgVesvQWdD21PLS1E+Yi0Vl
w/0TyXEB6lngHctVsYmK1uyjkbXwHZAbglDADP7uWGwKmxZmqUY15eX2CvxJ+pkK
pXEHOqsgH8JEyO7lgq4huqbTrdJfu7jOigoWBrhpp8tqdDUt03hvNMrop0FKXD7K
SqwUFkHeYLWRPGgnsG2uw9mD8y1zzUTYkTEuSncyb8uhUcqvDX+dze1kOtwcNqN0
O91hfVswQODFk8c8Nb1m0aZQxCDOclghlEGhqSJhYqN26vBKGekpEBXVsmJX4rXK
OtqaY+zGie/ZpB0kB29Xw0g1YTy36J3aMb/kYg30x/krnZQW21MXWDA9kT39sMVN
IKTMAMv6nzO45qKb79iTGzyX/i4HEXcM0LbLuOqjkw8PW3T/wLF7twkgqrM4cL7z
CZyLvGWlKd0n50A9/amP1JHS2K7xASmF6fClgdgjzL+wZGk66u6bfyJ5fWOM6vjT
7NaBaqvnG8ox0h9oZDC5H9h/U4xiEQvMbveBILWkQ1Z7E/pf2QbiK0UqoLvRHSvs
2zQ8y3LLAzlKw6eKfPqhAxXWjxp1H0bFLCP8VTv8pf/96wm9mb7yGh7tPqriTkZF
dL3p4Ys8+XKpmOsFCyinRnHp/ih/C/douzbCu2UT/WRIFuEGXZBktIVLrgnvuGJd
kIqk/HXeRo34bYWh67mXxYhmVCxyQgPhxU790pkQYTyxJHq5X3vpqH0Q/kWnrlEx
7ShQGhzi5fV7/ryN7RQdnhYuvnuZEMuKE+aL2AqYiVuqM7E7IuQ6hkq1L/afFMO2
FPbfHTK6SV8/v+/rGpR/nNDysdI0D4QylCrlLDOnMI/FTfJqpd9HSE7czQrGef3U
TAA/xyXTh7oQ3b6OEctdiY6S3OJckRR+mBVobUy39+ABedR2vp5QMATdr9uWxBcJ
Uzg4XQ874vcfT0BERsJiURTve3r+AQ2z//suLTou2wc7q4QH0C5fmZGGcd1bKUdF
vNYu6hXIWXIk2O9qGuAbg2CPAST2Pj3wi7jJSNKE7DDuXmx90VyP7UWHhuXObRsp
vWiyhIrKxNLmhxeDRFazv1/Ym+PL2kW0rmceU47B5cVY4YbgmhkL4J/5iFN2S3+L
+b1MvsOu/qGPWCND/LyTJbTZi/s2cOIvTj2NqdQ5HX/vGBWdjAK/jj1VPxoOsah2
CV0zg5Ec5olyZ9K5/yQF6iIgx/eDvOlDC1X6YuklvDIGAvoF0LXrhki3KIw2XvXx
xkW38kE8M/5qBORsARrfcDBf4PI1ZWhbfBcC/ClWQDMXdoxmg73y66YtIYwH1im/
AfGFky4fXlBwpICixgWsiouczXf/pql2kSV/ZrY0rN5qZ71oqxTHK2YZ/TxvdtTy
cJyqoUmWC+8U66HnFgcQO+lAdPws9JBJXtdSszrMUtGwd3gEDBEsezshEnouyeop
US03iRkpJNNlKH1QTNMrJ7Neb/dIlBIfulzCAgsYwHbqTzw8bhNcOcmY2si8N8bH
OlXXfbhK86kNqvDdP+xgyC5Lj7+TyFVOos9R8PXBNq/kgsxgIuWGltAMHf2JzWTM
Lccgvr9uA8DDw7mIenOKEs5Mj5QjlHe1XGW+8lMFJqmWkGgRBPeSorpwgppIZjDv
3IAKbxNtWTBINRm9LTIZCQ5JOx8Pe/KZ8WeQAe4yq9DqX1r5X56x9nZrVKjcjUe3
sujKdRrzB2uJeZP5vyBglDkcv92O6mbWKA5JIXV6Zo8OZkpHmjaObkkkl9k1gBEy
Sj2v+HN1cFO2x+HmicdFxR04Y4YIX62BQK1YhI8k1ZlGx0CZRhfBo9UmoJk7G6XR
zvXg0s8gGf/goFhXn+SbzvqNVJZgl9T00YkGYiFI5gnsF3/sB4y1enVPsDUh3229
eKltybshAy7tSbbDEAEl1URchzvwC9GMSZDbevHNd82xheL9XGh84MPFKxU0i/bD
rIL7UGyvzSO+inI2/larkhGrH/vJ5w5beSohRVNNjVLuJHb11GG1erGWYpw4F3qm
7e/vkTUaU9/EFd4T3hZ5xyGWhvpMYlKsTKzeDzJdQYd6tylINOYy5wvDXb1TNk1t
I5RdMyliv7KuItGIcDTcqfMhEyYKnquPgHqIq3Y9EsxEdRQaxGgfMVT5meVXdTlG
JXHY9v6us/qZ/xUYn4aBlGcEBg4aoLgb9vmL2vOt43ottdpdjLli5ZgGLPBa7EzZ
kWbIfgEnLLZW6epKTcxF11gbWbjZIOHUUaCXYFgReaQkksnwO4aPqyn6FJ/rQfrg
PGyxp/ee7+mHSFZKQYoLcZHhvI1UqaIiL+/jsj1hq4IqtBmPMtT3nBZP2Si+5YDp
Vh2U41Htpe34ACBh/g+xlMtfMaHkAIkkYySgaXSi99dqD3qdiu8Q+cs06qR2aVLo
MhQcu4FPIaKd2yIH0mZorxGoe/qF4fETbxuApRWQARE7fvUXidM44cuek0ncAKmv
ddWD41A/xoj/9tBUv/X3CC+lRmwrD6hdf5AzB00ASfKL78OzWBncbNtik96knVQt
IOl1+/MWs3dp+yGEFq8FlKOq9lW+ZPseBjllkNKpX52ttxebThx0rYF6mG9X85qm
K1P1UrExj36BiJk/LKZtx9WaDpAPi4BQ0Tg+voQ2nObxYF57AQChBtHyFD0oFMLR
vyGwSGJ5Yt4E0FtGG8JJhxPYwAn0NP1mJ4rhgAwQVcAMK7zbhzooWx9mTdFZ/vwm
LbB2KVbifzV6MUrPM4aFaBr3Tdk2736fibx+so8+EluPvwqGyGnIszR2dysOx4JF
LUClqvq1NcGmIxfSe84+PFMrZMPUNWzYYWJ32hdMNUE/GvdhGp91m7x882/BXvQs
0oCNpEqVO5f83xql/1peIBvQo49/VilB7lEBBZmtUkbuDAFJTzXAzhMyPHn4t1kS
PHk9+bGeM/+jh53n5iBmQJTIs1bUfNjMgkbF8oFKmedutjb1PV761Wg9yNj4HRPt
9cf72IQ16Z5El/E29F6PRKowiLj31Imw+/VXMXOR8C7jS0cEnjJztpI2bDzOWdhC
Y9amUFF/roBcAjnWY2hPZS3XHI/bL7/tRkMgU50pE3Z2FLoYTbqZScGKLfuNQsUA
z5erRZ7LxSDU+CtErSFNGHKY3IIPpn1caF7rtRcdHY1kLv6kCV9nq/5BQg4dXOlb
E5LK52F4Oi5aOKlkRr6ucFXKrwOQkf5IdRU/18zUOLINwyUFYLTI8rF/Evq+JjdQ
LFNVlV8dnEaFZqG4NSgIR8rqMksycx5pRibwrWgv/qiNvintd7cEX88ESkVWg1Qr
4YTR7gxKjf37ZlthbDJbQHFHt081MqLO492ZTgeehc6H3rkl6v8OKZEPv/l7+2s4
aThQJuvTHiJaOQVncvO/olcdCyBATH1LrS/k4T95Wdq0pWYmQ1lc78hgA7r6UcGs
fb3/NaBmukaLqe9FY9oulXLKAx8uFg5wqIGPDMnTdArM4hx0yxjBrmqOrWGgkkKl
O51BPXd29aiL/7WGGEfGjbU5M2hWoAwGd9ysfXlAmbdvcv8mZOgI4ALxsM/K4gUd
gX3lIOtX6LbfDaWU0jxMdablD4sE5gB/kNnSPkzslVMCwq4SnZc2tGc4jsJLpFs4
aj5hPAQW+s5wNxu5MFGKnpphJC12aRL3hPCApDFicoARxR6Tz9UHjEddQxwphyYi
Q7dLElSo5HMPQlOF3jusy9Uw2Cc1W9Y1IdF8sV6BCXNL7ePx/08jtMyz+lIVjwi0
/tWlV0xphECVzRWdOALwC4jANUnjNiyp8PrErkmgERRUCXG/beSJhCbFfHtmHMXS
0n+Dv7d4cZbQJpNM7dUxFLmPdHx6DFFUY1aKBTo5DVGuTsnLXYkYCY076w2fceSh
l1eDmzNhlJaVDKUALuYamw3EQ3VWwVejf68hVR5EEZMrT4E9PE/SHusVxQRTbXHx
o2yjuj10y6Jv26jM9BUcjGAASvUvqm6WtnNykDiZGbiu82BFjl2UcBAeRlfifYap
dLDW1PfiLwR0AAQ+avQInXIgmmyU0u4DIs9yZ1gq1uxMtx5mv7rqZJbRtWAJTdXZ
X8xjtVztpaX1LdKV6GgSuQdWQYhbBErUBzoj1XZJW3BkjhXyw4gDBgXEzYuaZObm
l8DQoYaPx58jD/vF87tLhusQNKQ3F9L5jSpkqGMWQwQHdgmy/pojvL+nhKi5HhCn
ap2gykpVqxYIOsu4zw/im3RZw4o2Svw1gurFkQppXUTZb4sgzOgIwW30/RfCezo6
CyhAsp0pkTVpEPKpyjFZfpLcdj4zg45qKNi8VFwytSovw1MsGgfHsmcKZ03pcCKI
TFJp4apkwTqqOYmmoPkzRwtTJnakgzT0FhkEQYJ2Ig+tkyq9E3rhP0qY3E70tuYn
ZNmBRpmef7UnqrQZ12qpnhuayO4L3AMptRzJZgmpaNJlgOYmnY4bDyYERNhDSJH8
RLndz/UOCaIB1YVZ+StiQ0S5pv7CR8NNjXqK9gewdhDfy3EZW+bLzt3xF8pyO1Ut
zsZOvB+Y7ILBfquSo9pfG/IO1uGGiIYxhMTE3VegEeWG8OcSZdG62dUEffikPNGU
R+2BNr+ZfFg54RjTzJxQIuo22yX4uUoUkf9RmLcnyueA96IRtUWTJXuf1Y+w4YYM
zBicX5t6RAmvJaOt+8aculkairL4lJ6qHxTm8/t30arVvYqg1Qhh90LPobNvBVXj
W/a6u04EhHykCU/juyHmH/jT9GUu1mMI7UfV7MrhnNvhGqkbClZ5x2GAIM01YIsV
cB1Fd1E9tc+cMQWSa1raNY7swrO20Tggof5WXr6vreDjg0nMMTPQld5JOwOwIoN/
7roqv4BmgnvTWNZ6QuitnQPkSDMw2GLI9nYwJ2qBjSgPX3Z8hADr7ufqorg3Pxkj
nAPxVMf2VQs8r7V6Uyiea5ohyVYAQti0j6UzceKrlXDMowK4UL3SD6mXi/gA8k3Z
hhPAuiy0UOD+lsRa9R9f3ujzvzj5ESuGT+E3+4f/MY+ucL+OXQ7ISoldF47iwn7c
Fsj1Ja4cPSFbayJFHuqRSFQhEjTlgDcgL5d2IkZZyFAFVVJMnmuNZFXe4aovet1Y
8/L+6ZlvEc2J23dyNleUniwRTM0s1I7mZ6nS2+FEN43mYFn4ddNmxlWMQI2uFWpI
CEamZsAeCCzS0LfbxaoaJnTIq3ECbkThpKYZrplVemW4+bipTILLTArE8EXB0qVI
PZQs88NRUzCd373D8e4WRtggdV/1Sf3Jl4Wy7ZKLqkFzD1R1GIDYebJVaYVvkZWE
BbjCBap4Zej9mixwUJjj/EHOzQQWMujEXIb9j75HBbQ1c+3nYsCN8aHjPqAXiH1F
c2AO4ZB3zM9nKLNsQGX8BZZt7MyokFJxkE1WFmncvyq4sL20SDElsUSICI/snSU2
w8U5FWk8/2EhQCzQ71nz4syMpgow7PeawKarQST8zqXBm5V57E7M+KNpjU7MFdeu
FpkDDiPAYAlgUHBhPodvHuZLCxlKXdWggf0ztspjFOK2megBhjTtDHrBOxOevGZY
8kvR8hAn5NKDKDbNSu7R/rJoypLQdb1oiE+crrHm0A+XTJHmGdLD+TxvVp+J3x4k
5F6SWnLrh63YDb42QdavdB+ukQX+KYmW1U5bYyzMmMilBm14ErgwX5E/0GX1hQhQ
7+nZM4FTNMLSMyZjWvDCLgtGDaQntke3KTZQ09sWTqnN0fq5WGn44TmrJaBAmsib
kMAygL81kJYZniMqCeJZJk42n4htJYfbpk4Mq0rMCG0zZbWLpCtt8iFI8eDb16l0
JWXaRzgI5XufZqINvQMvCbK4eHPaIkgOd+bKNQnTNyLLLS94OeWxnYjOiqs+RJVl
b+5Hb73q+CghDjJphwQJptv4WsApl3qYFzqytv9Ovi11fRwq7Kxh3pBhBE0jqiSb
BO405Gu1E/G20okJxgn/gBk72C4uZuBU0tS+eCU4BLek8SURfdKcea+V1hdfuj+0
64tHj7uVFDIy33t3rVN+y8deCnzsk8B99sVwRaSQu2oa+Y8ObOBAo1lstqjEEdH2
/hhBLLROu39YCJyqtuhZyxskV5fvnKwYDFHTtgBMDrefDosO+Pco74gRgjc6AD51
bYbJWke3FVNT402WxQWZ7B342Ct1EFVZ4T5oHWSxbSGgjtoAV2SnvW6qbM0qlfKg
ap2sOvF+BRY0g7f0RqKiySRFhymGanxsU/tlfxarI4QwkZn1kpFkOFaOv9qWOQzd
XrvMNFfQN1R5xRSi0oOl3DWrvyCfDdFQYCME/PNs66wQxVxJmd4kLUOF34B/V6QU
8P5y4lRXHsECyFmNARhlhPZyeV5LegmUxDXLtbb9tHzK77KpuHnZLTEVGgDd7vlT
TkRjvThG9fK4A4Rnxiqo3v9160S6lcrvCzuEu9H04nTGsAkb9vf3MBpfjgbMf28z
t6jeeGXKrXVOTolrhOr45mxbJEw9/UXggLnfkktbKZ1BLdgdyV1X3/6lRBAbeNgO
mXSroASkRVCAonn3O1a1RJEM8JjquhzmMusbURGv1E+ldQ8EYzQESFsocdRb8T4O
ik2VYrVnwEvUItYbV7Ud8UySgBJq025LphGNBFMp1AzMMrjcieaaN0vB2ult9rdb
5LujHPmsrLBaePBefge5A1EAj1ohdQmfNNFye7GLHrsRMg+eSBxyBx5Gc4Jexe2q
6LhwgI8MI8zmBbZGzzY4yg1ERAdPpLOF+Xd13aZM+srlHHRRge1kW4UuJsQtCIo3
ZXUbVDVlDdwW3+/26dI4eFADQGvJ72x0O1hsgOVuOWwJ7et0eOMxn8ergPT8NrxU
PlYHhZhk7Va7Qh0suUxJ3QTGKWXV43iBYo7aNxxLKsFYDsm8G63U3PvuTq3LPXss
cQbohe9DH/6bBHJVVijC08JRJCOAPXXz7yVzRmvV6uz0+SnUCPkpoqA/XrFbP7qC
ap8WabTz7B5cwuXu2Rj55+NF+UQntFd7e1H7w/Aaa5y7gYhH85pd7b3JTX8ZAJDU
tBgYXGnaG16adwGV/IkBOmpjBJ8gB7p1g2EN1qMpzRpjgAXrpFZNmaDEtayLpJ8D
tYeGmDcpy0xMBYABjJHffgnbEXMaIl/Fko7g476cFg0H2GgSN+/gjre/euVR1T73
Za5SU1FTB43LGD8CIFxFRUJ2x+L76rOWPuYl6jwzvO/WjAwwlIejclv6QzTJu/Ch
p7SBw0kDcgLLBSI1GFNZytIro8nrFEUEODiAd/A/rGWcDIIDya8nwDMvwoa5g0ba
ByXxDjHIz59+6GSxYc9sjfjkuaqzh86jQe6KpN7JJ8Vb7ROZH+kwsTn72n/WxMiJ
ImxOuueeI1ia7Lqg7uI8quaSli13SsxKMBzdLB9RyUoxkw0KazxscVXBJSXVe+o+
0MUAKFXkw0th7he00XjmgL+pUN8aIRLG/xMNXh8KQfbfTJ49OTvYmMynqABlhZrm
HX+l/QOtYQsMPvfNW6Rd9dxXTAZo4fs9QqgM8KNCSuagjDN9x5DOHv9AXdipd/Wn
gQD/lpdhTVyeNYFXNdSbJ1+gudj7l3C3t+xRE9nizn9oFKztr68t2Kiun0XuCePe
HvMiJYqZAcUhZkQEH6lgku5oszSXfr2WpOVDMY9rjYyMc3ov4U7FzsuOA0WOHrld
7QrQc1ACOBYepzGONuWGgkHKzuUFuKPjVVmB0CI6Rqy0B07TLSa7ef5G2wOJl16B
dvrME+8/89vmrgsFAGHmcQY0zAAU+tC2vQ1nMPjeQLs2ozrRyZnXWtRKSYErBBri
sl8zttbKiNUkYmdlmGqHDzYxRVtvNy2SOVuECIrXA7YOHRhPRO/qAe6gDlTY9f90
bSu3lGqkQ8UUeGzeQT62Pti/5Q1t9aFNjZrZrNMid56tzUBQq0NrG2fyvaj/p/NZ
trfyN3wdUGsKijUp58WatJzuCtE2LCVO55IqaBvn8aorgqk2sPykjUnJj8tDWJaz
Eu623aOEwXfwOXzUgicUBFoBN8T0f71edhAta95+6IWYw0Y1eWd1oC5UJOQrAGkg
lLDQvynHyks/fjsgP3f0q+xil0+c7DRxjsp5S6ybTtf9g5/AtU1rVL4Zki08HUrG
d16Xr2z8xjuBA2C2TcASys0kh+QZsZxkD5M74P62Lz+dnCO5028VxAT8biR/zyXd
MDhcw1oMt7OMOXYMsXDGHByw2Hprd7LfM/DA9A3wx7wr5k+Oyb/jn9iJ2OZH0Xv6
Ok5uROU8Vt4a62xwwkzLgGpg2CSHHpqjSNzIUkIFFywDotgTmtTYhRgXqPetopua
SuvmL41aBc+88fuUWyQBXg8kYsAIuGlKbTBh9pORV5sj44K5+XYUuAwkBysn1kZV
p9c/MTnk4vpuC0NHy/bV5NENqpIYpg+hElEWeA3eaiJCQ+EqzXWmIio6T1X0Kg1X
mccc/7JOiw8xny2h/waUuNuOjiQeyEsxa5fdqF1WeYj9gBFJdIy/P/Y4iMV3wxBz
yyVAAVTKaMCI0fNkD2Nl3XCAp+IHRiUb5hhYHTBsSoIEcUDP4yFHnNPGvkl+Lgya
LvxbauhuxwL1BMj52Up5KO6m6P8MWPrJnkKrEqRitUI0GE72r9GEge9nzuDYTWdH
998ei3vC3zwqzgCpQcN7ESneSoDZhY9y5OMVGdvo6d18tON+aZjifNAWdJOEBSAa
O6jQfOt4wKa1XPY9iHG+hsbPys0M9EiHSYTH59tdFiTJp50TU9Wx//NrXmhk+FAX
2Y9IUm73sgZ+5CRqEaACQtY6e0K9TNIeC2CU3S+h/y9FULLFtBDQKpmTPSvA4AX1
oeL2OhMq3e42lJS/btXA/0DEYBbt768s1KbdnE9h1C+LyDl1xsFs+W12Bm/K7q/e
umqTH9dMvFO3Cjaj4bCBMRfYsfzA3s3Hq/K+7WbvAueNoWC1Jfs2q0c73lBZVw8w
B6qvHP1LXLufoH9DLBcdUaL+hA6l5rqxZm3IgQaVNjeRz+IvmfX3RucV3+iGm3mP
3izlhCSxzGAofx5OXgM64bdNTZIocGD0NXqLDabvWC/1L7ajyrxdjnDZpa3wWByS
fRg7+ROif+bJrB8jeEFEie0Qmw5fvNfy06iJ+mPXAAJDAUwd/XR315D54qhJzebz
L1WxnYEeV2GyOmrM+r0zNFrzY2+CJD80G5Qhfdy+fEItwDLNSKmbkcmHUp8CecNC
gV8jsvPm7YDQjhOz65kRizwPtjg6Z9eTL5xrXCf98ScrrwcB5UzcLq62raBjgjZd
QAcoHKOqZg8MP+STpT/JHuOumeyfirI8ue4proSbVQQmyKrbRMvmcQzChEf21j+h
jl81V1k1/LLCJs4cFQ7KXxsKeuAgpb0sof9q4UtQ0bG7qMPvW6KS41E1k2/Apsfb
fZ9PQ0t52+tjY23F4TIToYNv/PKC45aTFX8dombTiakrmTkMBSM2Ms3Cl3MNZ8bu
matw7Z6s6EO84DtYDa6zNasmeeRQTgNuc+/KwjIHdFDdhEUkhOpIQvtuyoBtsy1U
weyIhlON5h++EGeJHQWLRKJmKYeKwOAecFzLPYP0SsnSbP6C0PcfFRtiuW0Sg1QY
jIq6U54lUaeUnJ/fQ6gYzU6GQEojUX0TnlkpcHRrUAZw0MaW/iLmQj6M5VX10pND
jlCxVPwgjfMMVZfOcDFSLz4VdGIidnIJnQNM3g0xtFAoHwy9pJKNpBSjmkDV4eFe
e27pIvd16tAQS/LaoA7IpPoivOpmvdHKKTmrwXXzPXWjflgyH/jGmrTyCsWs2zvl
mKyxH9EQ6TLO8CsokMKwc9Y168GgBeVh3cijxyhANO05GkUrL2fxtp6VR2G1x6aS
B07+kWjJAyEVRb7ACrldk/ulwIE8v8413vuaPCNL9EiUwgXobAlSkd6VGzrTs+TP
AeP6LdIaPSYgqIAoY7mvk4P4Cw8u4sOFk+ZMQg3iwVunTcwJIFAcxuRzAlTAiVNB
keeXYsm8EFvtdN8xRnYjx/Y2Io/z568epkQfEmaOMkn0he06NUM1TDXoWfq4yC/M
pzJd+AAiOiXmd33KzCNztHgHBYwPk1PH3ppGRRmc8/13k2Q1KzrGFnO0mCjX+EmN
AuJr+jR6QLoYiYWHYHaVSBmb/JeLg524irE/NcK3MAt2Bw17PtNO7D+MOz8Uyzs/
YbRHy2tViEGHAIfECBdi7nK3hb89PeV++XfgsxkUmt4B8z8jfsaVOsDoL17u9bwx
j06dHSoXVaIOIzcaVFkEcP8WtXp5vy3iIuVkINTpkxJN3WQ9mG+y+3ELdIwTXEZb
3KLAdiUhH+52F6qvIuoTisMwtDn/XKMtKklrwEiwNAyRJ+tGtT3EO13GlYmFeKqn
kz3jeHZLvIUXGsu0OvUoDIPt/TBEVKDz8aZMwvpvZvsl3Zj8Y6KQzVKGkzSGEIO3
8vvSE4pZQ3pc1rtXs2LbWGlhln7YNACVna8hvCteftSGKqGHVasbBM1M/tptRW3R
40tZ07VU+0vtA2kmfGcjUqeTJYJruqbaYT+XlspqKU9h/yQvjvEgDVlVwyaWT8Ef
5YyHND+x4nlMYjhCR23f5zhIZ6lOu1bYXOPmT++d6GNT2fsQ3usMV95/wHKV90aa
FBsL7GeDvI6oGmAkdrSqn3G0vjGuv++UoK0bTFJ7ecIHuwOAsV8hnasqHx4qM6W0
I4qMCDaro2UioEPg7e5iwU4I7QFHyPwBoteQldIx5IJs3N8amogzELOVDe03OqxG
fJshoxyk13He3k9uYMIJdgFfiDDIRL0KrGGmwn9EXzjlEMl9n7iSxPeWnVOCQzry
jl9bTiQsLn3P3e7B2/C3+KnDH5nACEm8KXnMyHzhnWKdPYt+JXZ41KVBImmDK49I
XiLhIQFKAinYhYExJi3lKQRAOfPfnl0lLA6OD7BbwWAvHfWFLrE3q9J3Yok8/Hqb
PSDOSUMO8OomKcdnte/Y6veKXOOfyqRLeIeMFQQrcxW9IvptrGZOB+mOC+KSAspt
T5o51fSk+z91KcurAJHTCwR19VfwpDmntXpoEpvWl4Esq9Z/55s+8BFdokFe+cge
X8ttHdMV8M8BUXVQvc7Gv46Cj/fJ8mV8ChWmQNn6+ay/hTWN/ae5FgbMiVD0eMHg
9VtbXm0tAmMuWPoxOncWBgMMyNWz6VOFeAwIdZs7EQ47/afTkYijrvw7FSctBKwS
4g62LScgNd2/hOWNCV7EWaccCw/9Rhhi/BH8ITaX5f5Ei8waRESIQF03i/5shGwX
qfvmshV7e2sBotuJ+rfG9pulRVcZ7n5rya6ZDdKGvt5Dg6Ci6Qlq3T6w8JSez8Xm
VFFidOYWIt6Y8iYr2QlCXs/MdxJzy/q28/E3yDcMsgtz1dSC+MYz3SBnfBhA/GSN
NdX/7A9V02gSGBLsY06EEM6bLCfRa5a7/vixUQzIciL0xzjbBn8X90kUlPAGfWPE
Ky6P5eTGC8hHyLJ7rt+MN3m+rjTifFFvmSW0pcK86yAKVQI+EWjG8Osw/hOfjmnp
F0U3mKwNy34Peq+MjNJBK/Tee1OR3MoEI/fN0Nsub+PVaPav0xrk5JTlp64IJxe4
mJ6cmTpUnGqdcGZHEqmU8rTUDLIRCxFcRXFzdD7GHb8X7DcieqRiVGZCMaUtOJlS
Kk9hLn2S1G1NdQSChb7PahhT6rKBJlaZe9eZegBgwFwjtsyj2ep5VzkXGux0uXuZ
jHh7p5IfXh1nw4WQRxUUBaHdhBdH3UFHFOzi2+w1sNL2jSxDrfwvnfNpY10S/PpM
aly4rVG2cCr29IGKfX88dQLnT9tCb2+Cyb8GkNDcKYkcYbs8LIIlpIEllJ2N+pr5
CeR0j4d97oEO7eXf3Y1wVPOLm3dEgM58I0LBhg8nsRMSA9ziq7GnKz1/u1VCPrcq
CQ190CIwDBydfaLL0XfQsaEZT3KBq4lv1oZgM+k89HDzjQIy6Sy0aOdwAHndW5kR
WMr3qTb3wEo1+axEF4AZYaXfAsEsI+4hJ5TstFxQlcbCBVgOdEQc2yCkWF6mYiIE
S7Rxe4Io9vV6Ei40kYF3x+ZpIEdPwAwTQS0QcWdWTZRRFuQC658cuAODbWmCE4cA
wHABG1sqPpxGjU6nwFlTQR0c7YVbjLCUM5M9NyOTJVii2UFaqLlPadTuUPE1aANk
hRhNTI3aB8QLUvaqPXNLe+QNtZP+SV9jraP1CUxnsDJogX7Blk9fuDouf2v3E1IB
5d6Tl2/xFFXi1CnQEAu0Gxp4l1WZ3n9EjRfWuS9jNTqZk/vmNGnpDQUbctf6qpMM
cVH2eErwe2Hig5DVwW3Z9+pc+5FoARvxykeWREdE7DcpPmww5vI0NgJ+yRJoBzSx
ObV1CP3vWGqYQWALvPUFNgnWt7AOz4iWiC+v2nXMc9k4LqpN0wMkpmKF2uytWyPc
6zdS69cTfzYN2dSZELuTSZ6+Elg96cBdqle8BRl4zuXNVHQ3AlKoaQhiP6CSc44Z
YgbQ6q1+B1oavzC0BsKxbTS+dZFaN27WdL81fE82BvkolOZFKT7QBv+kdjbG1FXY
llFpgBqlDZ+/6w5xYygkvQEx4O2/AwXoDHqk3OjvnA42lgINP10cDrq/qFMzWVfN
8qJlF91zCnwUY0R2yAGyYtT6MwXBokikXifWmE5fMR0CVfH1b+UEBf1nKqfef40U
k27gFHgmi9LZi4Ih+5za/spJ5axeUgOfg6xlso5bkxEtLSFPKMWpXuXgKTMrmThB
BEtWA3g6R1ZsIGyYLSZY8suLEY1AgEDn3IffcZUw0CJ0Ycye+AoT/WBcny72m17v
/K0i6QFAoIOz7nyBBiyn/426PuqVvcOR4xa3RZ2k5qiUDqgqZFnG1Mq/WeOize5l
rnTU52mIHh8ueBmnjYahtfJb2FzhZ6lmbeMAlsMomChaLm3vpp8rzML717whztPk
tUFsl6L82Z/di0HgGOlx5BfTuZqpFNA5Ic7ErOceGJ+esKjZp68/IusRWSPS9sHf
L/aZ+MnuxxzyBciczlqumMpPDiWkPInqzGbgtYnMtcp0G8mqJJ8XSOg7zxKwlM2Y
llAVbluV5TyjMo3SRSRNi6bDtYfwYXqs3Hw2mlBmnXmNIRtOFLrPA1f7BCRPVbsx
NgdOFhy0t8uIgOERk+8J1gbLuS0i/6Zt6RjzMaATT+wS+gpk4e/cSa6lg7AKvlgf
YCDnh+VsICTj5Rcy09wiDYcZEfzH4DNZneoqMJbYCrI57LDDFq+8I3anDH7mdySR
UxL79In97dtnhiMR1P3UdNT7NaCk/cdsvoZ8Mrf6dXKTQCgHAUxe28shmyowMUxh
mC2AssT8F1ahf/agJO5r3CfOTJFkEYhav05XG+fqskyBhhN982LPtiDtnr3JP799
a8WOfnNEKzJtnr1fsnNSOH6bt7d0aZoEgYRC/f2oWzNCAv+fYSJYcYeVbKhkRNTC
LiDgY+u1pKDSUWFU98wF5ToIswSxUw2USyqoCaEIc1hxDnrIfSXqftQiGQnmtAp+
fhtVvfulX6j5sxIZs03Zsd60EdkqS8bh5dypOSSDwjqTejLp8rd0ggiEj6KLKRVW
wl7uQcD/vIhpTFl3LivTZJnG5BwpU5pv6AUr3/Q8ixmn3pIvc5J+uEVGO96KGmQH
t9z3doaftVlSMomW729HqPfK4T64Kk2VdIJz+V7kRPyS3mFjiXZrcBFSboV2dOa2
6mWKxX06Vedh/BKFeq0e6rLag4Uko7qdLZ/ermE0+Oq+TSDACKDZiHhyGHUA9Wd/
v/ilOh7/3w2AIaDvuqX+N50C5X3R7hWQGTrfetkR0pnxr0opMnoP5yrVJXbNrraM
bltMIhugjC5qAfFfkN1mhAg5PfB7NnaFp4HmQ8vhQIIgcXBF0GkET8+6n3LwKU6E
0cA6B/Wsu+jCX7XQn74xc7CDK+/MdSbl3fWjDo6qnU/o1YMlf3FKs5psWkb0gJmC
AmQ+oZqwzH96AJDl1y2xmMSwXnw3eXQSZ/t7GHWnvZoOOEzjGAi/K5IUJyRB/L30
ka74OzAAd/FOvHle8cpo4XaxqayNb2hBLSykzPepRbfOgIhvhvun4LeyQkpfL64h
6QQfCbHGQVEtnTka2T+lyNJs3zg9B0jBsza2q71iovA9oL/GHhiBYu9ssWTx0lBU
TNNCSkym/s+YEwYLBFfJyl71cPXWZDW1nMxm6idq1/S4TbRM9gG5NX7H/RptAxtH
4gPlZmPLucAUEDeADQMMfdh3xjeywtqNK8fjm3Q8l73us6rmcEPTxmO7rREhrq0p
yzyNdfTq8FvZo9ah9anTbsNDVkfrn+RwtLLg0O9llXmDH6ZNWy6Y66NJYL3uHxP2
4aKblopkrPlblcJXpqb4KSkhF3eChvuEX7OeldbyifmQnb9aVrhSP1GNXNUwCJGP
x6GAv0niA5qVJZBeSVGjbzcqhLHqcq3OVGAQKkHpfoKfZkfu0cIZOEfAPCFJ+pVF
RPv9Rxnjq76JUZnHX3wK6KaM7i/zXez7D+QEGZ0pJTnBQH07Tl5yIDal8ffdbjm8
s5ysmqVvW+24bqCSYPRJo5NDJnPWSnZp63Kw9GwcsxoRa+/V4V2r/+KPEB08SOfB
pwAyFmyLly60l4Q+NftIWSnumJmwHyTD+2UF8rn6K1Hp/10vGF/n/1AbMPVFSI+T
gkqnvcvENZAwfXraKs5v2zA30wMQolAPzyhaLXf0fu7fTkmh0CzBv3EG/ls5Oz0E
GUO0HCFKlFi0FWawch7JWIigehDYLM5AlLkQDzSpwL0DUnb2yJlRIBbfrALHRTQK
nIx5t9LjA265goYBQMqGDnn85nJ7zZgbvEIWb8IjcaIKglGcmJMWpgxO5239nOlA
r5/LkZc6Y1uIV5/5BBd2fShulkJv4XVQE9VQw5pOaNyGzD5ZKgeyaTNxj3pUn9wY
6WvrbBZwiTDOd0LNfhgRwkKF9XKDE2EYFgaaXW+/oNTvXYmGXJ6OerHf+h5sky1s
btwACxEA8wYzhgK/qnvM6ITqYJu+Muob5+bzZm4PeDRPK73I5N5aWpXMgpmzmBi/
FlgLSGS9odMJR2do/UVV2gC0CsC4IS7aME9OjD5XkXzsiZ7HjCj/y5ZN7V09vg+z
qnL2PKeb2lWn0DkHzqNVcbZWrfNQxj1uUMXMWLnlJ1pXNI47y0xFhxsdcAUDcrmA
Y8o1UTmlGwH8Huh6bYUGLxl63o0pDBVoalgoznn+6UgUuDZYvpH9gyEm9IPIVHM8
tMC1Gb7CXV687PzgLZ8y1h6gv1JI3pX07o/zZtcx5fhsmtfrUGvme2fPwqxLXoPZ
QyXNuXeW2oqfMkID2WzzWWnFRzcNdnfONYrT53wlNqck1MBAql+DTYBhGpp9TQNx
D6muIR6sUL+KToQv8PAcHQPGxN0ibucpt1YLUo3yNizTO587V0qbTc0AeILGgcbD
Xh7DWr3ggfzoYhkUwNwTc09tYYcl492PsutciSk6PgWCfXEfWvc/Gi/V+e9HexVW
yAo2TfcKEs7bKGbyh25LQLHF6rsSBHyBAhZuxQZ1V/nF2UO2HXbTBeqEQg16UzNf
NOvW8tMNQFGTXagrw80QWimrWAHUUBVnSz1QSP8SwsLnZjmUpphNCFxr3kh2/VEL
XFqap0DvZW6O5LcREflS7b4f5u17SYOtv8Dis61ykgcXuiRBJfO3HgS2YFBxUOsn
VzpyD0yOkkNt4Me9hVAWvS08mpfwOvja70OAoqgonNNpS8EZUVL3McOzYVyNwTst
85Bpm0sJ2q/ZlBlO3b/bzCniA8iCIly1fXqLDBblYjxVaM7zgYs/hD/AbnEurjtD
Xbru6mnrAiw/ms2oT8QoYBbEZamqKxW/sNxAB5N7VgVWLBIz6V+9rnzy8TaNF7L8
fHLw2X47JK7QsvTA4FVUlXwbVTL+OS4ja2TSv4/fGLrZjhKPjGnv8ptZB53ON/UB
VspNo8aA69n8pkDAtoPS0YVVOW9yhAoSxhyH8Y2L6xbsnUtelEhXYI3gI8upfPiO
jb97/XEMhdm+QgMKe0mhdNgipBcvHwjqA6Dnq+f+lgFuheSzCmkaMlpSFvOVhMLZ
friiLbQVeYmoNE0vsTF9nSpjyLxRURJBP4iYAXll7FIuR9SEeWyhqI4N5QMX6Dgl
k+SzspCoXYBbrJ0URlTD74L5WUX5Fq1gHNDqNgmkSx4TY7peGXIjL+/9Vmdk/UnE
Ht5ZjsTsr4yT4kXu1IQuH/YWsce57+8g8xxvKA1n9ZVhF4W0UWmvhP05vSoMGI7a
u69czBmvSjoeg2Xe/fAiDIXWEGWKQ86Og7uaakKdWn8I6LL+0Kr5YOgDWUxTLUh3
xoPgu9sFUpp+lVVTXVguM698mhoG0amlwU+VKgAwgWgkNUDvnKqsNtnKsdB0ZJAA
rpplwcuDBJn9Y63ManN+Cn8WRIczkwnnrV386Xt8bpJKqKuF9xUZn6qZuaYVqqVJ
RuFmp2Rc+g3HRId9bFX+Q0qPiQBquo8CmJa9wP2/qbIyi+xA6R9jWqqLTltRo3MD
3w/R/LfNE2yrlMXuh938gi5acY41o+2jn4fp6ohvP4HLik26YhMDty9hCxPRBm/B
eAvY8tTQLxgHozKzgm9XxZeS81qzHL24/tWmBAX1vPINW0ZFAqJbgpzxPfhInL82
JtZFA+wLV+wrTcDPslWcJJhIWRbEV9bwh+3+O14Y4lnVohtpr3WexASoK2SOY1Ar
F6unuWYcQoB6v15QMC5U/rzSXbkWItTZB8biIXfCZPDIGuMu5spDhybux6XsuK55
R4AebkqduiWNmTQWtmkvVNGKnhgnTyiO6GGNLkktygRvDyV4Cta6lb0r+zFn/JmS
x5NnWurorzt/daY2TRZag01ubnawFzXPnEdWiF9OUMB11AlZ811MCaNRYru3MhoL
0XFuYNY6D5iecUrykY0LiNOPdM9NfLcgCY13iDMJki+eCFaLL4u4cWSzoBlQQB3z
sqFJba4zP5qg4jRhWXzJ6Hs9lH2AinyKtPBhSlZ7OZbQtBFGmPWUze/iPWvIsL3U
jfkBGD9iCigwOZvlM2wBV90GdkKAP/NF98b/cis1aWc9Y7hewf2t2/bWh8A49QoM
np7Yy0aCXKifFT7XJYJz4P1QcgrLxNdUkkAtMevLv9L+8DrA4UVmg4vVBXGyl7Su
XofeyOidpAgFdeLX/OMZ/sowSdtBfgpjQBnbvqMWmUmbhSuouQDj9Yii7QQUKtYJ
zNSpJhTdClUqaeHSthL8U3rk5fOxuKtHjhfx22gm2472MLrACwl81ZDgcSvtrhxa
3W1nd4g/EiAkQfHl/z7Mg9iMPDUhnR6ocMmLCiu6Ecs4+KnjsloJAFwaEY4xSmYE
FRt1kJGQhg8Th9m68nAzaoToIlEVG6s2+yaWWDRkVikVIZhMH7xvoK2fYqAjUIWQ
p5LHDfMKP92Z6OkvjKZCCMLWq+AcoDrSttIDVsxfoKl/EVUGgZkxz1kJjHvxv9rb
A1y1KI3SqDidGhP7tNUNH/SJ9UAD+60OEiI1VhWAO940kr3t3R2UDlm3iaGEp0Cw
lMbahVhh0ep4SYn08AAUhTiamR9XT4qf8ruOUHRFcfB6W4xHU8tljOZvNlW1MRUP
Im+Zjy9CVuSzllQMKgoSkVVxB9cp0ccECtzrc0GcEa8dWeQDTR4ArJKTOK0MtV0D
Wd7NOfLiena2uy4XJ4KRXLYzCHkFUh7hpSjBmUBxvZafM1673qAp13Owhg2IxZho
WRHs5EgnJGn8ij/kzDhpPYJcnMYu/tSfuOvtigKWGc7Q7J+RLmUz2QV+A24fo+f9
kmLbzWNdcCHwNHD935y4mc7KpyfAJd2A0TmfAfjXwFC+byk/v6NXOpPvO18wETX7
pp03BFQCAuOhr/tRNahh1dPfhTTjInOlN9Uowszk/iHGddhmn9aTbFDamFPh6muE
A7o7JE624zYHGMnxyWAQ3YGTMr1RjH2/HUprF/8k/ISiVFAdZe3h+7hhcBevSykE
wl90MsmteyTPOME9DRMKMz3FnpbYrzj3K+CV0YLsxpd2kJv1buysUgztGrWwMG1X
J5Pi+aEZnuaZ4OyEKfyK3LRq5th//b3W3Jygma4QIuds1mpVbybwuPGK/j660mVT
RGJLxGUH5bagsBnmoaibyrXTfmONyMDVQJkA9xEhkG03Ufhm/8RvpZUEPZFh+zB8
LVft35h2PbP/XPbqSii88dM2wfY2h/Vjl6VTRzLkH0w1aflbwFYhpeLFOG6CHWrd
tJCCtwADHcp52kf29lF9fh9JxaZpy2GqK+pvXtn7DsTt7AFXoh1AeQ2ExSNcErG7
6U+T1jw7RIeQ3/uj6QxAdQVHt6lP8xHxIepc2Hj++KNou366DKhu9fnfjcoto4DI
hb9/KivNDOI6Acq85CnnR5XLR1CZj55P5UXR99D9CVsJBIUfHgYzaq0G5I1HFRDk
hsHVX3K+ND7A7ycdTFB/XjiXNLHktnmaqC5SzAH8eMw9AFszlKQzLNEZslR/Cu+m
9nOkYYMWgEXjcFr77JmpDaXhM50NaWjUaTubaXf9jRf6h/2HLxARU/FwZlUA2veB
DHJ41tuxtBKrVOz1G3tdQqsOhgc8bdFvRlS8ZBCRqJe2/WHfn6H0W5jYR3buZAMJ
uEUjnMz9FgloH6TKq3pExgh6cym0GcnTk0nwbGgjfvG3VETKAOLoKvQP9A1vnfpi
bpGjIBCTxGqYJmBxMTjQ1dyMFI10rFQwWQTXyjyB7nYcJ9HaEJoH1h/zXbW/DZWJ
WxtuJhSwKk4lrF0tVL/xV3/Um343V/8l8atdpvVb2ry6uj6Fp7EtjYIySFH5dirA
Z9yk5V2fwVqiPjixbK4AQ9w/V4SAbHYADMpRxlpgQ5XryXL+uIJiiM0PKan41V92
hCSz7pln36iRdemfpmM60+Dm3ElzeYv1eDoM56761zsqHQ/MdKu80C25T51Qy1DA
Ili5jEr3XKcjLLvSMH19sEH8NkowoXCZPBLaN07Js4OhA4cHy4ZR7RbDc08Aa42P
31qtJjh0eLz+jOKpeRgAOmnttYAf54U5Q6pef1EwGMvBGQqv0lw9ST0kHk8lgGPy
9kZCcguipjozzdVh+5lIQBaPRomM7OvEyJfyT44XU3oKPZxIaUhLl2NW/6nDFxLp
qZSO9s5FEYsNJUm7nwlQ3Jbo4D7Oy6nNI6XCW2rpqusrLm0TZzbWIoEub5/7pTRe
G7wCDCXdBFp0xxkAY3gY+OMKGgi67sCeM9+GJMI2zSUr+n9gOZNKqZpro9Bp+Kou
nEOBC5JIYKARgNXiyxbuI9ag/GbyCxafi4hSOU9CROO4vpKQjhqvFpg67YVHKD7T
UoGyIJZjcRLMCQDrLcM71fOFhzUN7r/qtEMXZzgWIZxPYvVPRYJpoddbRU/R2f7u
4bdPE/esJqq1NDDWgw8FOnrkNFcgCxgVSecLZdPkk/QJN9mF6xX2APbAqrt+cCYZ
DHrstKaNw+2F8iNB0FhirgdNx41kll4wRmsEGF4MPCv7z+vPMNTOg25QWOp94s+L
2CRMoJD3Y0oYjNDWx0Ui+q6aEDomBMXeZFK8fGOiy5VUZEXWqxRg0/9l4HoXYeA7
Bv6ZxyR21QTqgW4c4uL9haTD9pu4CYNFXf4BvggYPheLFrj+HSG3mUB7iu8JtcUW
qXZdGV6rav7RSqnFyECJaiFd8KMh1vhCzJtUWmVIf6ngnnLlaUZoTqNTWdWJp6eB
Bjqa+zgYboi67EUm01i3EnH/8TD/5uJT0JCou1K+qbvVlcryIAQ2QGV0biL5CJlB
Og9OOVsuK0uizpbGTfS98MVycniOxNLHczMaxoN0fBc28TzOH1+8DzaCM6e5582F
gy0tsivdiLky/oCQl1kBb17SJuPuqP7ZjzektqiiBTyApb6WhQ+4H5+y5Mp65yCk
UYBCjEHzTcT2Q9OvDLAx5pJ6VONj+SlgmHZ5WZmchK+vx8gyPa7X35ZaN+8FyTgg
QEe9s2+6uP48CvDMUvdH6jbB4qa+0iyyAuHeHszQe7dv+8VqmF6v/Gc1X81DW6BH
0cbZQZSo/CTqh+OECgLuMSADcNP77/X5rGV4w5Ojk1P2vzcCapYhpqSdmunQM5em
spGvSmZ3W9983m2MUwHGQmv/1UZvDb7o7gUawatov90uzn9p2Mj0UyAMxKdrk9n8
oS33a3kll7vcfEZKvigilOEeursRgYyjDA8liWvGDcBbUgP018rs9t1ZQzX37Jgr
XADmXiwhLD+fcIYusFUak6Zk0x3aIyCaPYxUk92AR+g1gP3ApBAUeiQm2I99/rOc
VyY/ZDlNC4t0QzbYCESX4xIF+YROtJhcF6NT8ZAaBRkhDJvailfKWOoNtr1XRFNJ
5P0MOMfJvsHxQrBziqUxg371+wSRhFeQn4AJZJEaByslU0hYrsScTM9BSJVhnfMN
TaJrm1w7k1IQHMT8Q3cF5NhTeOQwEgfC2pnAl9i5TFOaePddFO2GgUneJaawUJQj
0suQ46GUfbZL0K1l6vhjj2KaKe/w8FXJUkqEpqcnyNjmNu+0KTUdrE+Xs70t254i
JD/B+l9pUpcGy+JuHjGYIhw97uwZjaIKwBjygg/BBXy3jjbyb8owSIdvsAHDBBil
COddU6GukKH4xecX/8+yNR/Y++bRf6dhQR8yBSxrIyxHsgY9bFDa3y99qUuafMFM
qeks0W89kofFw/xVw5a29xITT0KlBNElDalV7J3cAHPhRmTjD8YShGvkkjY0zqvv
Dmmn0WRIkLdHCvWFu8LvOKoKx91kHWmeAFea8XL/Y4Ityx1Iqzw/A7jXKkm8T+B4
uKjjVf88f0N99ZSH5TnOAFP+sWhmpbOhAyZeqgdRjo3hl+s7S7AjjZ+zhzyBvRwM
QaqZkPwJjJbCz9g5CCWfV83tbPcEUPTcihNzpLJAyP/NHBKZHKzMjWCQAicXhJCc
wF/3TA50T/48f7h6OqtTcgSZv/hhP32IlK/gUgyz8rm7IB4De2irTSRoed1xHQ2T
fB+LQ7lh9zugK1f+vMrJBDGd7m/ogvt6zTcMXq89pK27rBzLkaIQV735UAImw1Xz
DwFKixYgpW7yJHr21+phrPlSYdr5CTNV8YC6ObNgHc7CytivYZFe2OKySybg954l
JsrFgwJAG/qtw3giD9EQ1/MHgGY7DgLj7Y8W4VPrvJtA+S86bqKJ27ws/oTWo4Ma
BLWK70BVqWgfrElpMy9PgSCEPzJ0Ile9eoDxx54NabQistjQ4BYXEqy0bnasfynJ
gD2r2/F0I/KvTFiztLpOPfWzt8naSJ3uR6GeapF1uEQyyaOpbDfBOMcA7ukbwO7g
Bi8Ohqd6FCFitff65pkAAYPix0FTed4byj5HUPcUAi+bd6lohISDG3npSm8PcA4g
lF/OwhSLo2b1CiTq4pvN4B5Qd7L4+YZ3HKrr3ToOevN+YVK0LOZ6Pc2+0coU/9ZF
O4QvIkFJxWvmsyTUaSavyP6GLkZ88O25RXarzfYvayfwHmxF84S1zKmOlJiPaYb8
M0gHtP3pIrXMQZTO7cYdbQ/9Gz9s4jqyOF/jGNZeSlFXQ+MM3OfY10neK6axIBeV
zNojOV1ws0tyiIMobJsz/kA7pMlu3nLlX+6tywIOQfwkkd/WLRvQAGkRHmgF56ll
B1lZjtQClfvURK3kcsmAfgUFae7cJs61WpVtdnvnaFq0F+Zvv6/2PoG6VwhVCjKf
VLoFkk8ORDXy8IQr3HRD+zpMuEFoYv32HBQI8Bt5YefWqcmP0vCA8duxNt/aIUKu
ohUciZV/8nkMApvHU5fNg2gVknKb3T+eKXtVngUjP3KrVAB9XAAsSfm/ze0R2bG+
7f6WShHIJ3Sx2jfpr69S5RrGMohncUYa7Y2CkK+D6ZRqPkm9FXdELY9RDwkssmqT
wQ4E6QNjmGmUq+RbzTcXRAMheFhyx9VUyEvjT2p/WmoUUy2Xdrbu4jlzHcETPSF6
lY05KYD/syLmniFA7K1r+QMs8xkZQf6XpoJ+xEKND5ruiquxOsPZczJlvLl8Op5u
+TJXC2rd/gs99qg41KJuQhG6lXtPt+11kvNL/S72QUjw8uLBbMifSYo7KOTjNdGd
nZ7UuzUv0d/g04d7nDT9E3al2FY97tB3cLCGb7hSt2sInzxgYSSQBcas53pcgwti
SxqkXegevVGkfb1GotZKyPlBmlpfu0CMkqazyyfndnTtAjUHI1lslZwaW5ma9/AD
ff4HfMZEz30ebqS+MfwIO1mzdOzNCFrnRMIaaGNnBYaHnWTK0gfRAEp6kP7rcSfs
tc4ngyMjNBzLe3QmJ16shEiFmSFdbkDP6U7P/t+c4gadR6M/yeKjvOk1z2MIv6Bg
d0mRpObaeueUURzlJ1MLS7vHKTyUZera0U63sq6A48Q/WwHpuv+4zBhEUfbz0Kd3
w2cuVjz0w3MqefbWMNvoFCvln0ZVSN502KGpOQ7fDRZ6npMc1uhFPvzW4ZufEn4B
elCiyF2Ad0/dFqpfp+hKfI1STk7tlray17/k0SEEtUIkfx7y2QAU+DR4RIaQ7Bi/
HrBX/U8DJuDjD5SHVvaHDULi0iGCUDOrZ66HWpU9zIevjVNwIKNShTskdz3kCvn2
jubfNoK95jwqFcDbit96wviesEmElI7xxSgMPZnu2Se84eeCqGECahlr/BFXVwjt
bUvOrhTryK1m3HKaaPtJhcY3jmRNYiJs1z720WILApmgIx4uY0bZDzebqlRI5upy
PgJ5iXcOSAXa0cth7hJc10HX0bCN28QxqT3defzBII/VaO1wmUFjziVgp9v3/yNv
CyyVHN338KCr+isKrPqzUDu1FXi5en/mfZYwJ7dH1dggVkNd3a7YEtsNZytH0EjF
rvvDuSzaItEin/ijz1W+ICdZNUkl+38PCm1U8WYhy+nbk5ckwPJhWBbO8BJ9XBp1
bH329PQHf7QpcL1HxQ4EK6L0Xa+i8ZSQz2g9RHGhz9HNasfXxwWLOXeCHFc8xt1u
m19tsZihXxcGi4h3qZz1jF3/5U2Kv/Q2GCIqyBYe7flgm3Klxk0vhgMtKcdURtwa
5WyhHKfmAXJG5NqRqBmckP3vw0dHonGvqvrPYXJzqd9ritB3SAFs6aHiRQ2+Dc5w
ELiw3PQviNcBx5q9z945etKQDGm09Rv/l1fYUZugP+OdXc0+QJCUtnhgIdyujn6w
BXBFTLRC2ZWVC+0b1KcQEkq6T2D40jF/+VUBq7zEaZg7JZc/a+auCsjvaZLMawRt
Eylb9LJ9Qk3JfIAXBpZq+bjckg+1FJ0kJ0rBlcAYSibwTLoLVNHHyAmZc/jMyPGr
9ee5OJJSpISyDgB7DNdh37DFON06AE6X/dTJAolqJprFWJuK+N1j829OR029g0qK
FlePKAXhiLA4/h2NoPsxcVKQnOii7C3TC/fxcgJPFaspl4D2LCwLPBL30TqpL+5U
Gs49bPiM3+HC7eo3oyR4lslFqPVGl7mzoXMAxbrwFFIBf2DRRiGoUUo7mfB9idPE
EFb0+79a1hzuo5OJTgZhImERD+5Gipv8/bdRpT8QcdR8t8AyUzFHw3Jx2hxyLPhg
8zG+TJeL0gCONzhEKBP5kTMAMFXvnYv/fxU9BlUlVJQgYpxsa9+nGysLqn5fAYN/
rMvF5/AnHeZbT5w0basG0OsOd7Wg51Fp5g8HLzCLWPpuj13QG3ZzKDThWlsA+bWp
VoX0rERH4W8C8eV4Brj6jzQvLA+SQWGPGzNySfq9x3w5vom9NgX0iVA2mLbI7bcI
GRKyyLc6Q/wAu9pyaSCz2KC3SaD3azVDD7Rvs1Fyz7piECtS2DNzCO6l6h+Wc9WL
KcSHkt3jLrQIjBr3odWgK0FdzSJy3O3YXClvoCR35rB/SN4qcy69b5J16pQP/b03
smUJnsl3gVw2VmAoNE2q7ettKBNdKf7WHF7oGx1O3T3QGuWoYcFdxusPuSZt2iEv
WZ55bVl2Kn5qLE8wjlNA7YA2ZRf6G0Cruqp9Qu6uGygc9vrsixCBNzfvpOUQcWyi
YEe2K3iQTkprZDVw+LdWpNza7GMmz/yWJxHSLmeSN5ophfNW7LJPwnQICxS462FG
+Voywm/N3w2mAxVKzqaJ5aEQjJ19c2hrRia7O5brCS4QqPrwiMRlYZhrbIXKMDju
q+nXWc97tx2XlRs0Taq0fYFGpg1EMVh7RzFFlWBATMElY5PT/sRDEyptCcwImuBW
+WFEGag7ds+n/wEPgmcr1i4XvrMRj2PV8GGD3AorWBiAwewgsZqXIeQ2dp6O7ONG
5vaw3JqUhRpLenELe56FFOO0BaWcqydXPgFZexoYoH6zvNO7MDrgNnuBPxGQ4tcZ
dfpJnXtxbINx7P3Gxp/2KoNk0fY3quLcGoMd256DkPo1UlpvnXkrPo4wP9v78EMu
WbwwSW7DQUAQfUpFAIfwa1WsFKcX63G+1f1fLY2NxC4lklp8fSnUOT9VnBDc6OYx
F7KNOJvVb5eyQ2qB5sbMd65x7K5rAZgroFJljaSaEAnAGAfd2dSZazQZe3G+viFp
FqhRvAwTrasdMAlVsbE3dJb03UpxmeHuD3yL/y3LOX3TPa/oP3HQtvgOsF+TIbFi
GUCm/a+QhUYYl8w/i2Of4g5ZEd866LPPhwkh5qqCTW4uGa8EyL42gWpAE7mORT20
zAjAlt8SOl1HPJOIdEwnDSMTZ6W7MPwwoLtLpq+3ojahBKtrMlThFliyxDne7BCr
RiBtsQzPn9c5+Nenyxevyvd9RrtAORUJvbR0r7FDGKIR588ZXVRAwkJK6PNjK9Nn
P3q4Aie97CyigjXmSfaEedpgIqt6MYvOgSC3Y6C2f3cbX+gXMNrangR0zw7uD2ZA
3utz3NENzKig14NRepQHXiIQMSnFIRducRdtUmmSPROVDHSIOV63Hewpu5XBq7EN
Ef8oFWCQxyORn2PwKVAW+hMPRuklqt48HgdtP5ACVqSt5Az+U8Kgnbcy6cvSukRM
POB/culGVWLQ8LKoBQFVcEi/c6La50dVMO4khwSkAK2v2S+kgDqL8jIqw23dIMGG
IQ3LplMEKmFkyYNpdOP+uS3MBq3BrouTzpjP4ZyKeLZiocnW0br4RT1tvVn3s/qm
LiXXKplo9PWpD7aS4eaA7Lhn9dCcWZbp7RpiLLeEo4dJrOaDbKxrD3APTubGxWiR
AQRZVUtBbiQhNagCxFRb3uhCjWtMqQoXP6+aC8n6M/zKbDoC4feVjbS1XZhvQGzu
OzEWB3QKGgFr27vISvEuYAx/NfFop9kkGQFJC+oe7eivhnIuebpD2yklZ18b0j0m
41SckVOY1xOHElfnq2oBJezVawMP+lRoQ8tBgZYnY4kdkcS8Gv2ADwsDr6EV3FER
d3YT/4kz0wuXxgFtFMQjwECkHVCZFIm3xn+PCVYkvMUbOJAOOIk0bcz4oQAviXvp
d9gOa5pZ1PEO0ZP3wft7qjhMmL6xA8GavRXv9Q1lO4oXhNf+VHdXXrDQI24xFS14
KyQWFGg6Nj3ZRzj4tn8yl5mrvLAq0CmM0JVghB7BinTDUgwMNjZCuDOEZ2asvsM8
/3vLq8FX+5RtyJqX/VcDewg5hOekXTahRgz8FMX+PRP66te1sdPaKm8CP9JHzQeN
zJrCAl4P9xpcVmiibA6ErClLHy4FYV49pDH3XnGU4PwSRlq/9VcP0s11RtzbGJsn
+cNr05vgnXnj8SA1/byuqgSu745WjJ0B/GJPcrOBhBeZ3slY/tGByRh6FBMSCdDS
5m+dE2/qOUNRnsIG4VYcqFaZF8QXvKoKNhZY6vDy2gCMqMnSGnc+9rIFOSMeAeGz
XthfI7tJVuzFP0AGMfuX1sb96C2bEdyYh0EZzwL9zMDzrDgEYJk6y84kSt8obLHX
Qjx3TLzGTWRLcIrbsz1MEEBmEacorkXzLDn0z9xrgQJzG6zlEmhKA3eRxCpsyUWm
03+MN4UvaM6X5DqIsC6/7Xz04DITJzHhV2VjwLwJtGaB1AzO4ok4Fygou/GZe/Tv
MoIypmEA4Yxpb73Kjwv30Sd2KOVhRtfAJtBnBAQOO117C+QF+AjWo6rsjqpSG5ik
5Ss5FnI8Uu2gHz9GV6bjzz8yIR27iZ6lTjh3l5t0KFtwQN71MEQygm4M5NDduACo
KXa7thkxQYyQQV5MENWe80/jbzIyf2amUd+Re9jd3InEXc17FuASboAmHsBFOfwh
fdCIdFOR92rGEmN6RVXZHDfZJvfoUF2BYWpXWr3lRc9bnQY36XJg1XcP3JAVoVYT
uSwNzDRWpk+d4h7TTX5FljVyORuN0eV53EuwpG5h9YxknGEHVKL4Q6odqS5AyTEH
zTcL22fznM6Qt378gJsL5UStNTmY4vPFvh+5FibbwFthKkuyLyz01d5D+2PIa5eO
1mv/xEGBDBfRQOb1wCyZljEzZipZhImibLnjzEKqPzChE2qHAen+FJX0OqAaJ6Ab
91E3udXFKTJQfjgaEMvBPvtoxRbzLRScizeUjz4dGOvieFdwVa8xDRQ0dTLKFvwP
G0RAsQTziDvtJsLjyFjixQeMyCfnRoh3deEOc3vGs0DZwqJXU059q1BX+z8GnQh+
tvolO75EpDNYll4zsO+Lj8QQKsobwZWkdvuE+Qz0Jb16+M3jhJVVutyaDocq+QXP
8q+uoLglkd+XqMUbLatzfGiTxPbtbUHVzwMaxB5gUTl57etNpZJ6ec9DVEAdyuw7
4XDZ4OEjNOiLitst5vK6zrpPSm9QMGU+PDPqXN/ve8yDIT0Qqs29Umxc6bntoOpQ
NAbmxqAZV5Fok7jcxkavyhEi4HdrYnO7hj7jN49TdOYPi+R091suUFNqBTWelSwR
Z0RSw/bNJ2Z+ArUIDfwplUMvlIt4aW3JkFMg9+UaIAsNH+FrAdyx+pepK6/ubOV0
QIwR7lB2H5BUPNHiNX5CPclbHW8puLj9GhZgp1F01gGr8WI5LoPxOG8rzAJ4xi0W
58u7VS6obd2//BJacUBFeIQY22HHqrTlplV3rPmnppqkZkCfDSEKNdF7KHzRQ1RN
Z3ul8zSLMZ9VM0N4Z/i4v9fMW3ydIlIclkVvxIYorAIwVnMJBqjlpddr9Fthcb7u
h2Zg/ZeqyK9vFEQIWEQQBq3YibsvI1QjSR+zZFYTYTaNTdoxdRqwOWxfq2fGa4M2
x5a6GNLIQrY9h8Jw41uyNySoq5c8Gb78cdWXR+0CTh0FYEp+KEgw2McAKAe3zHRo
bV0+CRNV85NX/6+vktOnOKLXlwIhKaW4H6q+XDKANT0z/mcNbu+w70YxMokQLdY/
PSCPrHwt2gWvAs++i+pbe0XaxJEr42n/HuHKQJq3TSu48BvUg3hwNzA80P5zIh0/
W4tr+DoDavb1FpHJUnpiLe4Lbv5L+8LzSIqdPOSya2C1RvfgpzlbZF/eyL7q8TAR
n2SFTRgSmYzKFjuPQzIcakBj8ohuVBQDqX2bYRG9eULPOWAyEXwir1yilOoOAzYe
QCibI+6Ehz0e8goJhm1KmJthMuQPXPt59PO8Cs4Okc8pQBTbFurBqXDTMEybVHF4
2UpYQONEjLYwPNRZGza+mWE4JEvVdg85I9YLjZfBOR8hJi3KubBwG8UdDXOGwfcv
HwILRtr3JUcZR/L2ds1MwZV2cOLYw4eEVdXvBBsCIuatnAgDeayTUf79VVTPDBZx
NroXS821p0stjyAoXUQNriKt/kmXdOEmcbwRbFcNMvStJz/PiyZIXSbUPGPUSTOL
gzXk2mpZdGycXii3mw6kgMHyayjUU+mr/wSM7MfUzYrITbnxnQFrNcbBb/CsrZM9
TfVMDGMQlejnH5LuR7tdd5iXLgRJhhZC6wsCvwtPcx6pLdF7hwdi9HXZ3qK0QxOS
zEdenjduC+fkZ1nVgLeGGnhR/wYs972sUA6/t5EbsKcku4tT8iffhKDJYrRcbKhf
RTlWbCY9g2hEjNdl5Fq97MXBi3a17pJtuTSHNn/vSVuTVbzmpTEoJftmqPAGSfKV
UtJ9LicI9o4F9EAD7tI6NoZkBw2KhgLNbQ5A4AlburloyVeVk1cwllY2knzLO+SP
LFZr+7Uebm3CPCwKMuqVktJoM6XLEvy/gsRF582vZbVmCzs0AWRHofWwM4JtaYTl
ybAmhU3PLNf8OK7hvCdasv8dzWU0Sk1jncogzt4weKPKUg+/DzE71DLZIqL+9D/R
AWNqKfSS9CSHrk5WIlAklvscpJBLF4Kt6gCxvcrYCxzoY6uixd7dEZV7gZmR0avX
BzoZ3ETPNNzG7mIrBPJwcV6S8TDX5AAnG8eDyRlD0v2sfiwB8norqCSs9r6fpGK+
kbtEIzZorgimyZL0a7ZOhdxo9UE0HorL3q1O7nL6KvwrBSx8kbYKT9yOXY1sGeT2
DuoiRk5h5DL7W8CRTelSGkotDZ5sycNWlDQRORHXirg8k+W4tG3r3wD58iyhJioU
Yj0ltBV9uSuP9qOYovaq0FZ+IQFHIWoCeFGzmjlVe+ookOLocBCqdgUWVek32wsX
6/3q7Ups/djQ6g4IcU+ba94Eu1ppaRwOcAk2T8sAMcv9p4mQh06qGIiSespFVrUu
7UcwikCjtg3ik0EQWFPpWOH0BKk1RBif1/UVWGaLKWHVeYTYIf/K8XBRo0UlRy2M
s3y2/h36NFqsu3CbdnUK2PDb4gRH8PLSd6Q+BbMPFTTMha5kAg+B7mE2at5fmCuJ
u7PhYa2p+IAUUpVKto4NxVbMGh/6gY7Mg85s/Q4zvmkNR2oa/Otzo0p7kQXy1JkV
2Pal9yUzsVRTuII/STU+vGHkHWTFnjWpvysMsHUlXEE9Cn9N+p6D7EqCjWo2uj5F
RN9MZyhcfpbKR6oCYEEy/a0ZVC4ED04ADKbznwgf6kEFNfDUWxdE1P1wCFE0QO/4
vfnpCCYplsHuLyHivw7/APG3CLzmKtHd68ZMiq5B7hpBu/N38BMymAiCkfLm/JWZ
IHoX3a2bK61NuYDhRNVkoaMfI6is6lxaB0584pz0aT/AAep0U/CLQS0DBeTnjNf6
nPckfG9T1ZQcfBxioI75wjQINj94uw1I2AjBffS0+Q6MLpqT2ehornafEyWvxM5a
AmEfXHwFtAspinS21kKr1erA0v/uQC8MZ1U/oKN5Ix1QgMK6VjpVQmHw+RuGTztk
H+roxpovPI+hAjdFldgl+/3oh2hC0xzkYDPCqIdP8gelsJdG5j46sbdWQ6Ty7gdN
BkjKsBkntO/z3EUi9iOxLeBk7Ah1ZzyWNItE8jQCgfjObG67fZ9olpUFHNdaXzB1
H6Tg56RBHvCKzUNLm0avCsP+dN412FR0x3YQ/WMaJevcxCDQY/NE3drrjOR4rx2w
9Z1T+pwOzOHYgJktxO79vUvyAJ5+4BgwuC6Gf77TB/SpY1XYBO/4+yWAWXaGcA+b
fD2HVwJtCr+FQKqUmVXax53keQr37eVkvgyVdg4Ef3vz3Xordlo5wtsTatt9N30v
q9FHD0J5DLKohF5CRGqAJgsyfNvIZ8otGiWl5HGN0E6U32wF3yHRc2G2r8ohjwDj
vthsyDldE3Qi7evFj1+dbQ+LkVoP/w2PsRxY1hlAmyXPq1L04apOD0N4nw0tocQ7
2Qd3ZmibOt8HYKz5i++SbisjpwKQsLLsg8TqBGEuJI3KlHEUPBjAECFlaKxOjDDN
TpDZPVvD176xVYKGGFd49B406Q3yDA8M4plUZ/743IzJGkcctRue4pjTEGKFSI3g
ZPGxYHX2jXyY/EjlnUUUx3s8d3kByj/1VK3gNNWxWztATbo1Aw8trH7W1oAEM3rp
mjD4OiBuecSs6SeomVTZM0qtYFeQ0yiNCUsv9h4wa17ATIcfYss1e7B46oJFNVMi
ye0hkDjdeiBA+S6DL8zb8sqw4IxOIb5FOClRHxCMtjaWdj6qYnzepM+PvTMGKHYu
wIzU09lLzEAIipAuukjxAk/od9r5ixJG/Q/OZcxA1oUsgQH4SXKaOkTiS3GYtwAL
m+KiZD2tqVEA4TKS+znMVL9UCPf3J5xVO8XwIZ6psrRlRjFlI98TIwXWnjWlCL50
Koi7YwXjUf2ASv16V4WA+U0i9QvsILUrMSrAXInXbOZzL6G32svQiRG1ZLUDTdo3
5np/MobIRin4DcLzlso93mcMHayFDkmnPL97VC8tju0/j9NsL+sudsMeNFuqLUin
9mwJFECE32cHMTyncNUS7BIWGMAL52TUduJpj0MbTijtGCAGJGgNnMZERZZPkMMV
eeK7dW23q0+stiLeoshhgVkeKkOk+qUZUoRZAUBaevCe/2YPoRSmYi1WZfkctt1z
bclJhtk7FeZhik9QKVcIDClJ1J0nr1GRiiyHMwjYvxTpdFDRl9Gi7F4e1N9UN3sz
/kvGQ0k4rypR//CX8SjXE2E1aQF9mM1rjR8y/tpVBBvBDXEuz3SgRKawhJ9XLOOC
ISM0y93BgfChPSnAfjQFmRpDeK0DM0MA9W20LKSRcpNYsTuiIDN2UHz/w2DfNcBo
oGwWEL/y/w0CUZaDEHwZlXAGLvaXrEPZyxqNNAiTdH/clgo6USb/ZzLndP3P7nlM
SwEI8LJ8Z7Oenpjzrmd0oq2F9GuQuvyJL7E7Z08eccySPe/th9+IBQ3qpaVRICKA
bOjtdWZO6lcQiWkI4nEsL3NrzC3APjO7fJ8d+yXG7lSkDVAYpgEwEckxtOYgAAEK
jS1//eUH5LQ/CwOMVdaPjqimWbxdh7qJV5FY4HKDVwMjE4aCSV2PabfgVlL19h2R
qArjPOMuOWT5uJct0USuZjZY1bjAPFs5UmvHdXWFBUA5I5JAc0fi9w+ThvQk2323
ZeX22ck+bz7P2byPGCxsjdAADpfs2edlKhj1wGsiTaF++zn/dYW4rADnP/XyTSZV
2lRXbwXr8Mgw2T8Ufxt9JUI38adlle/03bJTYZd52X30F2Zy6jrnza7MU8ydSx26
AQZ562Rj7XfyKkxoBxTiDOhXx5BveRpjdKGfH5j/zegNFAPrTE4R3LNBk+9a8TKy
kIPUkFKumen+J6v9i9jgRAnMY+6FLSPn1zQWTQvcuQDWcqSo3r5Usvp89xl/ezE6
Qs2/RVPOeweHoZ3KoYv7kEjx3jZlP9FxMSAtH+6kzSzJ4hS8cIG7gOFGyCuat1rK
oHTeMBUxBgRTBDdo4JsZrvTJPhDf4O7mfXHMQeyeA/70GL+/CZ5X9p3DmbJcGZhk
Fs7HvPNkEfXQMe9g621VmfGnad0ldpSg7ERxmnhrcbSXVaGQuZ0dPyU9SoWCXzi2
/iAWtD64L3tvXkLz2BX7hnpF2e7/8lywo6/V1y6wQfH42VPjkR8yS+jHWWT39RcQ
h7J6O0MMC1PCA9tW8vLWOd14UVI4QYDCeNfYe5nfD2b4ycEDSij4bsRynWEpq8DW
Q3yp4E5+iZgPYv2abr/maVEQlCfi3Wu0GhzM951w9Uo91dUAiWIdt52+i0MGCmWn
VeXzl++eVpucoE/x8kNlJYLPGs78QJufanu2NLWAsCDQI9ia8jxd7+OaVOILr3jK
1LOy5p8Gk+vuOTUVj30W7xN9M1pi7C7hBaM+fyaTB3f3s2obGsKL3geioLPww2im
M7lKuW2o2hC21xbBh1OZ9PxtLCmItWIH9hgkTbg+cUW5Mf1YnmWWRukvSD8fpjJj
k5RK+QsDv7Uo0vFZK71Rd/LcxfNP485LrVsBfZO+2UCzET/qBuig76Rd8r/OyHYj
YS8Q52vL/1LNmHr1sb43UZdATdxBTORafMqaVzSCgm+cD41M8iXN6GMocEDKOGJV
R3/k9YIWbIa0s06XDqpZK8C+5ecl6sOt4gLfYtLUxIy35N95keMBNiPeK6dXXbce
dNYtCVMsHoeeCkwks3c+QPQYH73TOC4dy7SFHnNXBo6X5jP7/CTp6uIqbXqwKccH
9mebsbIY2zhztFoPuQ0wLBaYQWEucRyLubnasif/IeSNPeG4vu5ndOmOs7ZWDAL4
6PCVmq+9NrmtkTRq0/uyjQyBty8pFt6OsLQf5YKwpKn8N41vG8hwpRNSFHzuIcnT
B6xyA/WfMu0UxsnJ9kP5HShPSiiHqg8Wxcb4rY5pmjx11thAq6v1UOKyz1DcwCaL
zUZkE7sTUWaGI/XC4tEXHZc9NkeOgjAf7fa0UwfccyGfb6avgmhHkCj7+1lUZVdZ
S4vVelnHo5pjIrXJzI0rk3BUe3sKid+7n9et75+JK8KRQBLkzPIjIJkF3h5TFiNk
cM59Zg3JMOIxSCmHC4KMnlxq/fJT/cpt2zet3+3euCVyTJi2JYe++cdQNOekiokO
tPGgNPiPXUSDtEDLos4+eO2OGYCdloh6e2l+XiiFDt/7isqGg94exh7J7gaZ2YuY
+bchOA825F8YHZ0C/4z3Ou1ZXPzLvXJ/KblYhLTKW4CvnT8eCVLG98aCq3LPz6jS
9RfaymrNIXIjT74qVdYuep1qCLObMwfySXkJAXb6yrBxXe2hHZDdb6lQwly8rSMC
qXBtmCAtp16eIC99kufZdnQzb5H4YocCqrN3FkCCjarMVbyvqpuZF8kZY+BAlAW5
3WydJKUoS9cbrTLkd8DjuKe4pyIwxtoWX8sGzSuccMvb0eUbB1qQCL1X9y70kKgi
ec+beUAjkg0dcQ0uop/G7gEL7zu5xQ9mcSZ8wOdVkAQVvVKyvYGaxsw9hz4E0n9e
tjDgyRZXPGDW4KiRY2Ir7f/FB3/r5+Y6uej6iKuPBsCR1/hpnsD3OtE2N8HN8KaW
6DlpdHIXB+IcR19GIUfanH/jEmtbF5UN8FVI8nS99Gbw7bHbekhOOW73exffUdM+
AtOJvxEmoqRMfyd5x+YaMepAGOyiwxuzWMxCI6UfpyG1Dz67O+i8mXTVSWMgYj67
N7yZ9SCr9WS4zKEiGyWVoe2zCVkEiPrSCQ6QnRS1VY7M9Ysn4RxWOb/Af/DD/9em
hZMI0eS78btCj7rkUAh5U7Lk74StYEcMJIDyk408CDp4YW9FDCWWPLDxLJl/Iw4l
6m/qKSsaGWxcepp0UA0eIiktMWvqFNdae0nzW6ghsREuWDW/EJo7zPIDcaQSgej0
9h5v3Ed0xW/vGyZXIgsRfGsd4lQHQEaE8WoSQBwTye+y4Lk6pfq/Dhq3AfbrRYFg
xlYTYxrTIvNbv2C+/KnawBuuFbiLQRE/nPoX2yDqnx3e0PaJirmQhsT99y2cvluM
hG5BnWYHREL4llTPwFrn5vzucsb9m1OTsWmP1wbUrIIUVXSA80QgMzhfGnyXY187
QTlDsGgq5/LMI/x01EG2sJzNv9aMEeHH/VHVUpGC1l9+pfAjsFyoWyNiQpzAmZtf
p+2ULOA7OVVnXcHzjWxfPFqy747c04rDk9N3rcklysuL21pS8lyYMB/SWISmMfVK
MmkCkK1os9IwkjT+fBDnWjFEGkJ/fX9xYIftAKlMVRuixE04b0XWD2m2JrnM2hNc
kWv42Wp7y+DZ7dJ5ySgYPqm5bQsqMTF2/z2r9uW2ULCugEuP5VziINCZ+919LXU8
nP++5qhMH4ECnwe/NbDwNRZDtS7GMjCf7cQExbcGZQkma2doubeRICa7Ha8f1hd+
1J7UGbZjDl+xbQhSiUB19kcYqv/iFuOf4xUfrD1zpbEjjRN/zch3qPXCrmDRmC5s
yiCTE4vxFXQitQnzL6tRT6GmZrWazqQMIZXDTFfjKsNP2uuml/F/wyNKF0czCVNZ
ZG1Q8V+aKiC6BtpKUKniCOxhpOanN0VIVpTLFwFxV0kwhNFg8D18LSFSEHO3qYtT
1lX5kyNpTX7WT07FKH/0rVkoTKwUv1KwXNN+ufwIXPuy/OPyVC5nEOkTR5BGAKOf
hUJVHWRmaGcvZ32Kt62At4lSKsqo+I4s5fKz5UrYNyeSb5ErJDgLjcA9BEQFCt/n
kURod0dk9ECZVPT3FqCyKYJDciz90CQbH4Sj6kpxdaM87O8joY4oypxMIyA/Y15g
bFdPDOehoxeMtc0htMM6hd4S6kO8SUThPeCk5zmGZKI//xOpCsNobqU727eCcAjU
jQGBU5fQGLt5VfNQr85fovoMut0O4H/fKGiqufYbqs0+gjalS6pSvJ6k6Wh3RgX0
RMYil4eU5ONvbz7iGEg2gdPlnO55XLyfhrfQerEEHJ0VZwuVSJevEGOtmY2o+vQ/
Pl6+dNrt76aJ6rL2F4K/ruQe947JDgPm+eruwFJhZB2DDLe17Tr/HChkGtlpNXP3
pheuOZ5O1Vik5r+HK3NkJl+wL2g8oFRFexZTSlK6jwnrc4w1sZMFfHbLJQpdCK+2
QaMFgJFGjCDariM6bQrOjUrl6DJqj/yymA+HobgUfLpGB/jDvJNkwrbq8IQeSecy
AO4X2hhKgA7ZZ6/KJ9MfptSnq9YXhEZ1P9pKtq1jxZ/j9kyMoKiJ3TX6/OgXupK+
QCB2MpSSLJG4SdGsnU+R6mahCvSpgmqCZCYVi5UxeO6ANKgqEuZxjCyDtzfLBKPc
nlWG4Nzs/Rxwahwkn5chaRVZZoRQqWAtLF9KDV8Ny594zayCQ8lawWnGmxeM1Cvs
hrvAEKRAmzDLi84uzgynyqZRFEzCOXJZIxDI66aCSFDiZ45KsRffNMeGbdG+SdJz
bdPXUMC3m1PlVbu5jGtiU4Zqte9m4k8T33gyKROMFlBrVrMZZn/BqwcfnpKNFks7
sld8+FplVSSHmeJ2lHcbQIteFIHwZ0okUkbJhB2CkFkMARPd/uBqBD3P3hacWEBq
1JdzlGAhuHAyqXpYF0jjTBMUV5/6n5Jxv1YQHncowa//1USLmLhooDmr3M5GIgGM
aGA72FfRO3XPdIRw/+rF2ZgYG9MOZa67DzffDjDk/8VzV2whk/DC0byydrWg/qo6
tWm4j7rJxgDMfJ3uVoGGXUjQ7l8THzFbwPmSQNfBbo3VJJNKaYM6rQwUkeaim8vg
WEsp4mJwIMbEky+Yh5KDb3vdTowXEIXJzJhgZHW98kx8uoVG0S+Xzz9Z8mms8C1j
xQinPHg5o58IE/6AkAECW6BP/vJkJt2cBoS/YFs+yLGsfDnMKzA/xRHpUyWSAcy5
kc5ES9NkjLvwB8+eDqcFrl6kq/YE0T83mHPie+JXXa9V0uKVf3X+VeWK90yaBDoM
wI/stwuAxpObJ2cdcv2Wv6Cw4KyxUTRgfglTT1F8hBkl6MoM5nxsCA1bhhOv41w2
hbJPObleqzBrPt0a5t6frQpSsgEokQYfiNP29+SPgYqB3iNCZkuRg8YQ4azCWYFd
WDGBt46qbMMWw5kdmoyZLM/M4+/Bui2JAXN7o+ZVugYGEU2iwWftXFuWlF1kcBW9
2XAKsKpNURiG1OjK2xy9KQm5j0KTBo8SMQ9b+vQuyrZXPUVRD7n3IWEkguTEAAf1
wjkoZHdWUwaX2OEYWhpGibx6R6NT9eCU1p8glzOlk8YFf6zXyHneLDNy+Gyc418z
6mjmaBp10ZVXMDX3xVGdF7BiHLuDZKko6Ra4QQ8yoQemusHGLo654bAYR6L0psxb
ca+cUfigDNSm+J6TH1h1WYH8O/sjJPI/h+k3qUKeSPK4yAvQCu1o/s81EPWEhHgq
1uLa+kfqzy6gRdLhSIH6NUNrl0o6Ky2SOl/Z5RG8947HX359TdgsFbqwiX44msDV
yqnEWSsPdWCe//9Uhz54bKaqm9wB+BFMqZKNo0zs+NbWZd9xBluwMGM6iohNd4pP
whL4aB8JCtx0T3cm87qaWRw7Zn0NvrQXcWErBUwgojuFfiSGkEthT1cA1vOyL9/+
0gMX/9ebgE0PERv4VikAegWRGaOHyRpvIIc64A9UFz6VMi5B66Uwje5ETnGl+Tgn
vVRycOEc9GuFkzaAWzV8EaY0Fs+ADLGGl/yBvLlKIUz0WiPSM+5lQfq1a3YPHkqX
RToSLLGNFIzRDyYGiEeewKwQPvxbx3vJr/it3X4yW3TzG517CG+BFR8Ev/Rr/duK
CHboW/dIlK4+UW9qqPjTC+Q370Ipl76aPjF9fpD5xQGRTiXPiiR7ttR/1TTdM0yj
4WZ7QxOw0wUraJQnRyTrTaWLU/BVcZ/TvAqnjYrT3xriqgx+09zllnbi8gQVAAfl
JpPyfAYiK1+VtRLiLc86BQiP3VhrvK6E2ftaAJr5aWQCeYKVTef07aiOIzs+Rsdc
pqBvSGjTDSkDZQqrWVoqU+1Pu3y5RnDVEzqABHU8fjI6AzV31hiNWdKKa3BGQL7k
yNKHoKhagZghDBr4V+vWYVlcs/ska3bRgGAyVmPYUo3Rb/m/mi5JrJ7OiRMjvrNW
Ps9ipozCPqZc7gAD7JKGu4ZJ75x3u+bjMwf4aKw//NdFP7hlEkjURPkkOOw2TWeR
4NwY0UYWv7O3DSlHxXwXF+7RlI9TsFNY+pxV/t6BwblimWgBnSjyRMCJ49QJOuRK
oU8d7zAeKKjfLGNLmFkb5RkALZZ+e0X3hgjah7Fq80dpggZNostYn5O9EVOoSjR4
2vhHRa6HI9pOgoK9HzSVZH5yQV5xEg/Be/YjkofdHC+FLz1WN1wMzuzRUViwEGUE
1QHpoD4UKSBtLednvUK7BSVG/ER+94iMbHEBmQUaiR6X8uG87+zQbsMRzEIo2Nbg
WMb+ZehNydxWFUG/ZC87ffE5sApRhzef1JzgFJxGgQ1KvxvK8Wy7i5MKpw/DBacO
FT0nB+AQm658ZXATsM+EDSkjGnPtIVSZ0cM20Hlew90WmEnVE7WOAdb+kxPYmvVZ
BLOeUAKmCcVN6lBaGmeA2fcPPe15Rvqyid3mWPvl4VLY/dSBpjVmMWNTSOPXL6Jc
NGWJFkPCOMf1fvoYIMOqHMYUt4WTnle+5+aPPMesl9TbvvefVV2r2JADwEPfHaE1
lxKVN/vrn73W9CrDtLThV/P1w4fjZGb4ChcQXdmJvOU5pMJK+N+jVrKKiJx8kQAC
wu0dspA21TTTrm8IOJkCW2Wnq7TWQnX3rjQcWrBahVchwya5j7NJoOIGPDpBIiEK
aVVGSpabmF3jXx8Vv8M1cSPt3FYfOtNHGJZSLNpoyA+6sR+XUlPuPe7FET78GtaJ
ztWLPfH7tRSZzgXODkfwzLEJKBNt9eSocJzVE9f6jty7W+9JaPqaRATRdusaaEHB
RbR7kS9OaxYBrW0IVd8lBQAonk7ehUvoKGK2EBop/nPWmNvmEunf/b8mDQmtUQXP
V3wVUX4zTuraFc69A0X5jxt5ifUytlhy5A1ICdeIiE7eBeL9mdXiHtpFDnZIHvmE
v8tYIC9EdYByhTb0aOVAgH90AHpJV7QF2L1I/QDUkq/UyS4Dj/mkxoZ+0rz9/CSt
7NLBgTFxE1uqQUxA9leAGUWX8l19hNipQrHQ+D/M7qKvv2bhom26uWTRqRCw6Rst
hT2E1/LdQ0q0lwDP6ARHffvuCxUMp4PTBeNRWiAzhzQZWW+3Ie5WAh2nXNx21F9R
XnPXaOAx0OuED8CL9r65hrV9/bgRE/ohMuEBMj6jb6U2ySXfAyExP/+g6CUgsPZO
PrmoX2xR97N+uhYaWOMtrm02y4adKd4ZP3RUP8lpdWtrJtegU+Wi/vA50hRpnKaf
rzw/SzZ51KUXq4wm01+Zct45u/q3N/SnrVbEakZaJEHe4855ZW6RVZT1W0UwLiAU
figuYNlqcfV8xe1uWC3/IrY7N0DITk0H3YINGZCDegHk0ctbOy+iyF9gCSejIXg5
Ls/gnszhVaargN2LiwGlM8b1oK6EaemJTMAdzDCcZP3kZpzu0lwMB4AS7ETIHc/v
Uphoy4uTSh2mxKCY6qw+GYGMzK0kJ7JwjQ5FWb8aAnqYip0SD+Jyt7fxAc44/ca1
aS9DSK9ujRnhwGjNZQbY1l1GgYQeJ6VPrss8ewf/6s+RJpuZqdJfR36soJYKH+Kl
hmSAT4tlO+VPw4IcribYbRHblibXBr54qtpV9nuXI3v0R68f+i3DTiYi3R9f7Dva
B8jQwjhG/valltb9h3w4f57dSgr0TL3f0gJX6gQAfUirwUxVtMtoEDTHmnLi21JC
twUP5g9srDxgBEeovROLvch05yTs1emnkfPCsv0XoNhUtaMZj+C5VzOl9jW5LDzn
h/Z1oCKGLF1vKS3Z5RxrwerXLc0LPzpDTyUAVZqqwIUYIBciAV40eBR0DXhxYMqw
B1kwhttsEgIvd7w98HF4VP9kHjeUaH0VB8z9Q+pBQohhk5zGJtwP1iLkkhPVqXAz
iU3eJVlTqDb/ZU4ABvkpKUzhCNv1+6088hB4vfvT0YdjoVn4zGrFBBGN/qa9UYYS
nfMji9vFeXP3TVMkYJqUpDetKOlVDIt8ZRZtyJOgkDJctnXBhAzvEEBmDfIprOlr
HGA8ozL2FHhbwrzdNPRq+63mTf3oEIiOZ/Ex9CrvkNRdxcg4AV6dd7VlrL0IwaLG
HClCaeuygQO88exdgvJxGJbqxCl7udAHYEBNoYPkom4f1BT3rnwLZalmzGWW5P8l
ZjYIw3JSN+rilCF/0htd8nFKUjqy9xXK1Lz7bUZWYJ/cw5Wmf0vIGYOlCFzCKVih
NLa05f8MrXGNtXRCNyJcmnIE7Pmau9JR+Wyxxc4o7yGAhm4TyhjjaoQv/Aleiw8r
ywGKq1AB+BK1ltATO8x/tjP1USmMvOUeqY4qUAtdeWR+/K5GGpAOVISQK2ZJ0sPK
olimyhBN3ciw/zpgt+mgdQcuaWl1thmo3TM8EBRjR2AjhihzeAQaakhx5OLG0UJO
mxwv2v1J7vfogpjxuWmyRjd6kQHmaT7w9axSUcK/ySHoSCNWVjhPZd9twc4hyawC
eJzj9FDN74MZein2huvMZ1pDTl+8UaiD0T3LZVAcR+sPDIRNIYwXrYresLdlY4ns
DHJonU5tppCFqrRVERZdys/ia6fVRYXMXaBAZ0sfFnEy54+8F2eI5XpxlSREgT8b
XNUOHEKm3N7gKiXDlyM8c0UVQadc/hKG4BTVWWzJOq+W/Yxb9JyMpgEF3ph2IIEV
kNPMPt2GdAHN/vSpkEG0IavNjv+neEPMaSEhKmP6iE1ImkmYPriNzyuvdAhj/atb
8YLN6s7I8kzdxbcLpt7C4O40lQcUvrOzmISlnSorQi+QLtI308FfuiDNNMoorppv
EERnKR2LZ0sNPnwPkDKcizx8DksYYxJcrSVNF3WCIXJ2GBZEoPCVTuakL7PTq+UL
nmBX6pFhc1tACyS7rOMLFWvZMUpBUJyNisppVkQmALAZDLfpR96rjajkXRd9FEle
nHhrSR3TuwX6qNZvnKeaQG3AN9B+ifpPvmqeEVR3VdWL1JlVjAdfuPWDGW4GfWrl
eSdDA33/Lr2Wagnkz2FjPHLosAqcwe9/8N23gC8U4mMpZ3KaztGVC0OVAZSe4XMB
Rvq674+IIfAmXE0as5KFkFnqEW7lk3pPI9UNnwgCQhGyAUqQX8BARRSXJAkw4dBH
gzXWglGDR3asVDjZUzkYHdky4WYNYtJYIHVLMS8hDR75KDe8zDg5UeH+Naxfeobd
pjYQt2LfXTog00YdG+PN3kuf04QW6R9+Te6wbN49R4kV6W9A77y/3i8FQ95I0Luu
FPhI5Ykol3+qQtWnxAZXZA5UJmZFlchjKPa876b+dFpRXkyg7+qukImTMFMI8xcZ
F828RziZploMydpX8MxiFWFEqerHnNgyorpQhbKDxhdUAhTYQIbHY7MQlIf8Zt2B
AIz1m1MfqvxQnadI+lF+M4roMkKdE7O7buEuKumXc3c1QLCzqVuJbR7/soQs/E5d
mPXKDOET/2s+3cCou1lUGI5SvDyI0VSngM4J7P4uVg474UfsgDEJXQLXSbdSuQOO
XADllHeNJxhf09D0bdhoyF3ruuVjC0NV1jtyw60txMMhKCzFMc8PfH/7bOG4NjCY
IRMc7CnJIQN7kCiT5LR2nlOkKQnfVstLH96tmiVMtT8vNihrHFl0WNuLUsK4nYBS
uiKLSx8aYlfQcyc5QBXEMgP2v4cwdKoZ5kNH5PWQYCJ+aGWK0ztEjQfXtqsk+bWU
IprUozMXobyo/ZAYCcOsrab7ktHsiuBo3KRRXlORuFv6cdUw7U4iOq5Ie7VPxd03
4iwQS0Lk9LBsXLFuVD/TUZrp2mmTDcYK6qgIR6EzRw+i2q8pEWJI7btbezyyxpLt
Odo89yTPoDDD+Q9iKCYlQjdYgbPZNg8SJoZ+7g8jmN5H3ZUfBuO+6niP073Lu3lD
PwjLZ9pbyjESYAWmEyh21Z5u52701/NA9BQ8lCzzLII72Dfh5F9dYGxi1sEmIban
ulwySHglZ0DkY0kAbWBrRyGlJT7eSb6INy605IBJ20TgG9jXDqsmzxL+Y2N2Q7wZ
cIutmbI4sW2R0LDzN2eG9NXVf8JUzg6C1na0tc8RTsWD+PpX43yOavdiI4UT9N7s
96iBlx0iU28Q7N3JulMqZFSVoLn395x/HiycPhiulq4xB9jwhxvRfTlOQoe60LEg
SaPK27AZN6sa9vzxv/Xh+MPBPdjrqAFzoymtYN9h2c6pl0bl4J3kG+GeG7q7z63E
v6uVOCafWP3ja+cBHrjRhQ7TFPpwp63M9WU3HIAS+Qyl8PxpFCgOwJslRDROjf7T
gG5yF4AViamVO31hzBpqiZhpsO7m8KRbxndMLD/lvZ68oITrlD+s/f1KS+M3wvih
aZc4+hCfOhJzc+DZ5DDhG9ayKMDM/QEdLzYViXD2YUteTsP1H4LmL77sy64AkJu8
CLXmfr6ELm/utYLNwfZZuE1ZWzGZFEtP1Uz2kPuCBmQc/Z5r4WJwuds5L3f7gT0U
zxB5o08URyi2xrkOBi6QAW63I7ImLv1UtLi1FSpvNjMosQhvVJkOXL3RQ6e/lh06
IiloKDnlfFsbsnHrETEGe50ywF1cJaYDkb1iyH1RmDnxVQ43Zw59JsLYRr8hFwEF
vx00/Yty4NaoznZjv9HTCpsY8Vk6zhA1t+QxA0KzI0op/DISfaJgpGhl5kvKCYR9
fXiKgI3rnVs/ARMtoQxS6QTQZqGroDBYKVyOWT40HuWaqZefdt0x+TXq3Hy8pcOV
4eCekyjoOFCPgZQ9kgoMU7KbVef2caHNLzmahBmXQ+7SxIFiYndbbLulZWrHco4/
oUkX22UN+/t463rA7FI9G32NaGECKLe2f4vvHEqCmc7cus5GLDvBbci7jArEo8MJ
MmQNidrSA5Q7K8s1ZriBwFV93RxipqB6kJrG2bONs+fPD2z3Vz0u/G6x9pm+ZHDG
jyPCBEd91Rsw09CchAJV32jUx5ZRw01PX13e7Jx7gJbg8U9PFbpomW60C5UaASEC
wyyDsiZWtptFh5YP1hIVFwOYgYrNrjl07FRFZLpvv4+WmWHCpQZ3Bf1RPDndGjC1
opwB3OUo4UWXBzeYD8lD6gRfYTPlGlIyK643T83yGARIgrFggjkH2OvGCmE4dFEl
Urw3+HGpNgIx7z6Il4qqINtHJ9pUJ2s2JQCywgp3YFri0egy1swjCMPiXNF4iYJA
ttA0yqPSFtdejmfIWFUE6G6UHxoZ3mcXgDAVfzMQ6rLFzlm77zTyL/7kI/J1pwNq
njYWXs8bRjAMV8gq37vURBzaPTuTDFEN3T8sv3IrTUzSy1OVPfrZKFND3OUcwsf+
Vl3Y6z/RhxVY/JCgwxhpYyIR1yrLhA+fvujZUZ4QTdg601CxDqncVP3o0X5GO8B2
NfGdIEPLfuS0i3B4zc37RfxQ+leOriR4llCeDFYZ0eaHjciG5gNXQj8djMTw69cW
g7wHRhVXtSLS1/qwA+EPhuqOeD9d7aTjQr1QRXSLR3UWYnViN8eIGkpr/XoqVdJ5
gSgZDKOmrQFM+v7GrrZJnXN1FbqnC/CJ7QcmaXwLqJkAm9os4cm6s2CTWyFmuWHB
IdUi8RlFQSfLKn9sqTzUSYiJvxjQw3hQhF83Vhgoe81ov9tl73eonMKNwW4Einc/
uz5TkaKIEHbnYArB58F3+ftMxHE3BaJd+YE2g4Jwezmgv0bQRHantQbkIEYlEO+y
AoH9Ilqh3pZCz5d8QKCs3TzYV3jGnjLKDKRjJzGjqy5fBZzZj+anBdjRSF6vJLMK
1vjSTRLBoSHNQ66xDb2w8g6zDmR30NT2DCAcqRnZe20R65zEoxLSPR7P6IiJrZss
X1Aq9+jFUa86hBe3pxIiQ6Odl9nDWKZvYyOZh7gCzjk22W09Qfk7yl5KVKjiZukd
yJuPA6PZYiqQLEobmgkLvDtGsRX5/Q5LJc2860Viy4DyTemJgH8bKueXooIvCChX
i+rO9wQATym1wH90iTFTtXJUX9cLW0qeXmSeKjuBCRmtdOb/hYPtu9HuCKXbLjS2
mzDJAui01IcLvaRI7PAymmhyZBTy1YoyRP6wQZvfp/BedLrfdgFx5yCueElP3VRe
Nb4+EzQL/wsf+M4tF5zxMoFV4m55HvlD9cCWnRERs7SrMeZIaUjakkMQobG3aZ4p
JX4vMzhy6q+1oQStOIGH1zIml02EbuXS0o6XJlFYWPBJOmWjsSQ79Uq4CQ2DBROd
drXTzmvaXhdGOZ62qx9275ekC1TLVACN+QIRDAiwLsrMATVarYVvWKA6OXYNKJEs
VAm8XL/VGezeBDGCKe204as8G29UcygOCi74YqZdoiyCEmDLkEQgSePXfFhHWIRi
zkfvxG//lkqICPF5anoHfaRSpVpVyiz/IqHTKHG/N+LnzfdOkFNZ2llrZfzZp/mz
N5/5B912csjHXX7LGRPl/Uv8ukMxQxhNpq2Dgc3eQu0Vp5VenYGSlfByO+Oj4OW5
jc80APBnZV+Gwreuo3GPiUsFdy/qcDSxrYVLWELSkgqJDK6rA4ncQymd/RiEb4cp
BaRb1ybcdmB8F/L0HEOWyYyrZWhiaH7rL1W8X+uf4EAoCtV389ajvnW/LqWg0Pzn
8JzQ/zg+FNaO21dO9UWeGY7M5S/zAcD+VPEEaj0aoOtZbAX3kRgu5+EQJqxSxCVK
EN6ccEJIrc/c37nhqqJfm+fJen+E2K0Fb0iQpuItHlLfXSj30GbDzge2veQhFleP
JxzznksK6TdJ6aV1T50oMoxTDX2HdMWUf/yhTJesv3IHpzCDeEnqV0bUHlDc+8Rf
qUMF3SLqIHM1WEGbfPH/frqK6piJEZWIQIWD6MH11b9vHPZOns76ldKvzdcfPJeE
YwKTLbvvyil+x/QVXCh/6x9dVTKzHNakDoGBrzt7YlT6Qr2RIyZ/MPaxepq6vxH/
gUKAuCbD6HQ+9uOFe0Hz3hX4b8a6NIL5rE7NpywjO/YWWrTlyK84jyAZfwKKG/n5
4QowFl739h6LSsM7wQNuok8E7cCidJsMnv4O6y4p/T5l+/wBG6Q1zxy3aVOGJIsz
TmJz2f8FS9KpXvVvjdJx++cBQhdXkTvKbPnuhHgBO9ZFaTPGcBi8G6+/B+jIShd8
h0AJtW6IXkSbTvT3e2AHnWhl6XgMRIXhTB0IhEpvmByJRf3MS7e5zog7zBYBjdMd
m6vJrjhQG3r1Lh/6NTWwneU2CaQEvn6RbdybqHQyR8Gcr2tFzp07X5u+Qi40Ujg1
qxxiIvSHdEISpVip8GDUJx5v7tac+41cTRsAeXk5YR6mOjpY0VJOI9L+toGZK8IY
l1S9b2vclOK4iMNAKFpg+XV85xS/et96NYa/8K/pEUpgmrz3GfW1Ai9vU+kT+a2j
0VLqFsuv0AKxxPHkZW1hWkxUIw2F4AofssJxAe9o/Tp2/ihjWwmKLwMW1j64Modz
whHVISmVcecNI5k5a9WjQBSlksaStUO/jLAB5XcOaO0nFE6W5zyMAuXvvLOIXGMK
tyYPg9RV7N21JWKCl5nl/W5tgZbAelrTyS66HMK0p98ApYbloMtwhRuCPwAo5Vrn
u8cgoEEUqRsbt0rtR+RpJi+G9k397nH4z7M5tkgvtBtDxwoc+w4JiXf7rxXtxrFB
mbpCafsWiF4V4d5Uog2EpVbEewaBIfQ0qET+l9rFHstKlFWRKGhJfzqa80OvTaNq
hpBjcbQ3H/cGYeK61Yo34eX7yet4N8y/iVAVOYeeh4lOfp403tOoKl8kzbD7ntbU
tn3wO2Ds5yr34tdWQCF6gZJ2ebWurAJO2M0COfWLXk7z84g/QxggsQtuvxt8EBmr
tJt9tyuYeffxjzX5PBZLssgT9MgZg7rgB04yxxRrGHkW02mEyF2xyYq7eHxDklL0
GZNtuFzWo0El0n8mWfB9Nhq6ezxlM+8epGgqOBeTPPmrh0gbUBtEbh2gHBpx7TDG
K3pXpY203+YYC77Q4hSMxHKZbDySPt/gnU3/+oE6e7ae8m6IA6rV/kKKbYy0RYp5
m7bEbkWiksIUQn6N+7B/OnhJSOyZihWwK5IcnkkE/lZO/RO1RiaoqF9OAJC3nBuW
Tw12nN8eyE1NZnI2cRtrsyHKbLk3nQQSHA4959AZu6TRajq10LCIbSVIACt/zoeX
uBa4Stm1VkFJ13KXGEB8ytYPF+j+wJ3g190mj9sBudCEmykf6hJ+tQLvMfnjlvnX
xqG5AnQoBPZircUa7zS9Dk3xb49Zkc32p6WB2q5h+fp+TP5jGYjMGFydUo1z97M3
IO7x2bzaZGMVRqkPp0SbdHpFh3a7nYc6ZPzOFJNhkLjE2pLLo84lMp7fwtiJoBT7
kdae0/TGbgN8VUY7sr1+q+LB7rYrAteuBg0EWligZJNRypzoEVzGgL18UmfTxFIW
GfjDaqQ4GS13zUEF6QwS1sd4dOhyPDC+Lyueg+jYmtRHw7JmMKN/BfaKxNFyGfQG
WmvrxxkUH7QVHr+7Qv4QiuSmqJMuRBr05e7A3sPNy2zODTSUttQbIKYZcvSU4Kub
kon9uth1Rs/97kOyctA94/Uj1iCgUPRZm8FVLNS3SG72Dee01pIiUQu01oZPku+6
SYPBbqnEaT6Am9eubWixZMhhNXmXeBf4x4zXqbr7PTWzRQRXLg0Rlp0oDUTtODk+
vYUMfo96QWihQeZJzJO8ejQeZiKWgwfXlZoIZjF/UHxZvbvbxV2ByIglDYe0Zu/J
N0hQR/YfVJNgCXIzsQSZgZhBWOKZmV0beRoq4mzQDXtuAYpBnu6SNG/TptP7DrQX
H9kwLO/3wsTEH8mgwFNO92ewQkM7WsoeXJgvtKAfR5fUIYN6+7on3HAh7L2rF10S
QAfwXBeFwgSx8HBYXmTD1dOL/YHKSclZdEbznYj9b4oYSEE4CJ1eN0aPUpeOGviN
ryzDo3RY/UqHlovzI4V2PlOnDKZzn/oFeRW6n9c0xsv/AcK+OqSuC7pEDWIdh6Ii
TA12PZgpytA7N2KlIBRptvjLp9vULRiXZ+Ha/rI8cfeGI4VfOLDFYDoQaOR8+l9a
RmowX/bktFJYyI5VZkqWxYioJWKGRFfnAYEARRGJ20DpiDuFrzbHKoRaCeUJoBAZ
qiEiFdC81yK1nTXxCO5DniqVV03qTlUZEt7037bGvnZeL/JSVPn/rAARPXeYkiiB
yls+YaTYoJYVId/h7T1YxXV7jVDyGsL7PuePCTnf0tTyOgIonCuFG4beVE1NjlBH
kCStFbIPJkdNtAjnjE2p6BYSrlri3udvH8fk8QXAXbl6h0OEaba+yx0L8MdGknXb
0RNo41K/o0Ea5ynrKEKjTUScNiCJvMaMfLdzogNy7tvsXUgMLa7lpr0lCQdnhcjr
7zrmwkWEuS4qht4awWMgD/90aLDtwSAKHng2MKbgVhfJutmyV7oyyIkxl3hh7S6G
UaXji6nAn344yzPvqfO+GZAH4JNYc8cTdCNc66BBCnQTiNULu9t100cQ4ZjgX4rz
VhsMEKUBX4RfVd0YMTnXJVGlhZumrfjZdIax6oQwGPqqOuCDn45+ABEe2/PBl9cq
6YT66cYqe1NFu6HWCHEXsy4IqKFe/aMVz5Ya1/p4vPt2q0Vab3nkswJWDWsfRmEF
zWhcvJY5QqZ9OgrUbFmsYSW+cLrKM6uRqkqV2tkim7oBUEJ+Ypn+QGH5t04Kpsde
oKOgUIdkrt5W30simq55BBq7qdnqRqXDCdSCacKL9Bi2D2Q6N6BOS2Fh+++P1gto
uTIdiUYMdF9+Ey+XuWbvP52wGWt8wHVkJp2i28hUMnT+MKrfOVxrQRf97dFd24EQ
nwHQtq9e4JtdyvLWskQnk2EPwAxwToXzAIs1vOHxuN/ek28Ohlwp0y653TSaCVcN
s5mLExokf6S9MR0g93EO36ifCUnXWuMYs66AwVaX7XFBnw3i1qxWmN/D36+npDYv
G8HozTogq9LF7Oha508jS5BCp5r6gRJn26phxCeOFiF6mVKfzS3iyP3/Hgmd9ODM
iLxjGKlwg8a5wK5GSZWQEsdozL9gcJzKRQZkg2C6lBTg8PY/RSuNgrFw3ZmSSbqL
aoXk/2Y3rJQlBEHofaAwrp4dZYkWN3U9VphR7grgo6emUXlEgKumi2X0RC7NJEDy
BTZfIXX7agsLcMf7KPTIC+jwzc5yzdRfkLcho4g6/BnunsJ3POn7i4luEEh18kHh
a5VhVNLykBbYKUwYzHoSG7uKSKZofFHY0tYkFTWasUbDQwl2+TD3zJGk2qgsR3NE
Q01SqXgkDocO4O9r7Uatlp+5CGBeUp5+EsraN8G3oW3cxWxYiHGwVFA/WU5wDH14
PrQhUQjoXeDt5sV75hupdM5ErdpO4+Hm9cSBNQKupOl5UEgizMzgIWgCpJiQ4CID
NbXgC0daPdJ0tFapzMrrnjYtuocKvknKAzpkOFeY0UXN/wTUzjSpyCQRLNAUQxng
Pl9X5YgVraR7fMwzhjO0Uo6TbyZXaY+bmFkTK3o/3SY7SwD3H7a3xA+9e0kzstYt
x6sqbenMlS0fiNed8YoQ9DvF84CVD3Xx5ZVZ8yBYM+LTPEuoxVbWi1YK6pMT/vvA
AVkStuAw7TvsXWfUAvZFlmOgF0lA7K60cqBIIo71A8mBgKRP4rlHGvgVGv3aCpVT
BMVXL5e58Blgi3eRfbREu7vZNLcqBwycYag5Bc1wkzRQfHb4VJpfDgs72+1X4qZB
I8uIv5Lo5eH4E4kh7ZHLizi9RoY6Mq6Szd6JrUBjWY2MmddzWPSnr81pwmJ6tDxI
12tb9BxLYdAnS3uRBZ0bGk23L6HwCwXMZJmQOrh41iX8UXyJ0s2JCVAOLdg1szxl
bjURgQ1P1PQN6+JJXwW6y/afPk4DKScvebNPcwHuyI/+oy7cjqRrzyM6ykWaFjM2
ZWQFU6VP4xG3SEJJshR71z0jp5D0K6mp5EPkRRshIwZsnAVZn+Imh9fxXQ+HGOro
NRyEEpF3D706rFGCpJtzw7JF1IWJebZ8UQasnlkWX716Lyf5+KoxX603nzgDD4/8
kkFjxQchmiUozPWLbSoQCWEeY48zbbrlPrh3XcW2DTbKywPNlyQuIf0pLvhUJ7H8
jKDkOApkwvx38PG6FlQEU2vrnRBEWlgkQfRW5YfYVs4ZFQGMnYfsIWf4Kv7u3mYu
f4abf0z+ym95fuRSuSn8VxIDqPSjJvdSdDBlcL1nELBXLgdcBXH0g2JTmbDmIk2X
jGO8x6CVneqOrFz7wPD+/jKuf+Pu835C5TnwDM+HaUaaDjNF3IB8y+71lOMOdgH/
DEjT0ojaWGrMeMXADLAhw6mgJd9WN7Cjg4jKyeu8tgliN9Dp60uzLGfxlpC9HxNi
doERWD0xDzDb96YNv4t6T/vUnIfkEs445Bd5dFgESjwBp7JKmfbqQzXcO+P2yqFc
99JSbKsbi67j6IjQhxeSZsxZv5B8qp9nARY463JYk1W26oEV+c5Pa8tA6OQai+HJ
ebqYGk8f7R7Oqpd6v7ZruuZOA5rsmcjOSXO3dVc2rrlqC0RcTtHpEOps9vulfcOe
0ZFrJ8nPEHJk8aJa2/mfyWssTkIkjhfchUgo1ueQR1KuNcyGgH0bjtiRh068S9Ip
OVcJ53+565jlcFYFcSSpi7cUhN8ebabQJ16yHzr+91ISOTR9+tr1/m6ulwXzbAiG
RVi9wNwqFOmkH8RTqYP9MdyAjj44bMXqZamcSbgua7dP84TuHJW08yIhVywvB2LP
3eq8E2NIDMBmeFfF2V8vxFkH/ba2QfkT2iikCmCtnSXIAqtugekBuugsRIE3oBni
LgZr0rghd7EWeXlSwoZpG3M66ad6rtCuXixR4dVhw1SEWHqOFszZ5YS8WRlXF63j
KmRVHoZl/qGVStOtIFrmfZTA4DVqO2fiLuyBxzZTJJubdqVwPqcksmsreKo1UyoH
9CnDegEJFAN+5u8wk+hzLbiLBSPGfXNCqwHDS6eaQjTo30p5N2oxJ4JZaqie34dS
KvsiOnbR5QfC9dGq+W3ldNgUYc/cZXJ5wiWr6Gxyu1hCofrzxrUYxeyPh/46w5Ix
QfypOVeFSssaTReZctL0dpj54GWmztWlJvq4nykrwd3ac4VD93G7tqH53zIwLGSc
5JBjJsOnZ/NUZUbcfJJWc3gZfPRCFonZBvQ1UnPEekldSOkIaFAA1YzF9U1pPBAz
Y6SsR//5z0mOnHFRYCVxSViWURmGJbq571STow3FGQEcJyvSzNw4/iW7P0FHC12O
j32aPlVTkSVKr7/YpsdzPLyXA0GmGuNHb1Rjo+UU+zWXavK/lASjwjsy21jZYFxR
TaBkLaY8acEXsKhXOB1MZqnhBaUKCM6s+YpJuAlheBvOz0FsxdpCORGPKvrHClzI
RrUUI0FUpuIWb5tWCS0jveU5B/DNdAibyTa+eM7JziQJa2FGz6pYuPBE7akpT4Nn
kdH+nOIGUIiPn54CrGaCOh9CLaQdiTRHCB6hEfDBmbXXcocXFfqiAnwrm6iaUtGs
9uvEDwxGAG100ARGp25oI2DCUvz7XFCX6wby+GHd7GjTG3j0wXX4H+7Kza8hsfO7
VQs35+St7Vycac8kOw/X9rmGsq9JFSjaktwjmHjuU6pp6Qskd3/jXVwD4OWZTf7x
zw8nr3qMEz0BJUznnzHTHcQ5NB903W7b2/R5U/J73NYHkXKaEsc5bHud3MsKX+Ox
kAZLw/E9Fww2kjeIA00JlzPbzPAo9A55L877Vy7Qqts6tW0n/7c6Ul7B5IJnPRZ7
2vIzjlRotucmwPW4uVYzfwOMH7aEUiFDrjAx7e9Za57qQ+7IYXgtvd/UUfHX2qgG
IvvWvqi550b/GpiBSCl8Q0+rOCs8VP5xC4C86ZcldL1LGwcp7Wo3X2L6NC2G/y2h
LZpme6TwJ5XupSrPSFt60RE4P09lk0InNU77N+0CaPX5DDXW9IBnMP+tKbH/C3fv
npJGwRU9Su3OgVIY7ifIN/Fw/VyncDcwy1HRx2znB3Qgkk4fi3fMD4RNct5g4I0m
3ZRIdo/yoiCoJBDN5rWab6VunmHN9xnAkH/VZfsggSY/F9ar6SN84fSeL/G+VbmK
G2EyzrmgmG+Qrz/lVQWUnnGCg+qZLpy/WA8DKBZvd5ofzstFBRxLlSUL9e7kQzzh
w8ZkHJiAkYWXUXh6D2BUAIlkHVoBxY/s5xSLcvWSDc6OEMwyfLPo+Tbu+t5A8fcj
xIF9VmIrWBFwChLd6UBWf8xa3JZDFqZ5cQ4QcnavJalzARdapgyB85dlHay3HreD
vHbBY26uXFB+YB/vPz5wszGTZGNN1pJ/Sz/vl6j/0rBXf6WH4j2qKYojQ78W7CzV
0h3t8bFB+S85+Z1tlG6JZ84CeSz0f99EF0xQqeinM7yNJNDawWtQgHXux/LP6kVx
rlK8Klu3g1+D1Liugb/3fseIP6hkTDJYIV3aPHfGyPBC1iZLdnMwSV8T7UrO+jLR
aVNlhrZ899vsJyH+KIxe34R3EWbYVg6CvGxq3wtjTvuf84dwuQZHDpNs6+YRjuzk
Yv53AojafV+Gddq0C0+HL82yBBuf0ChSO2uVardmMeFgCha/+NyrRtqw6I9xOrn5
ig/qBYc0/pQ0cHjjSRxSGvPGxGv3WnTJitptjIrm9EujOo61LA8njeiz9jsvBXmG
Xyn1PIu+TIIH9mEUaV/ej243dhKusZ5JXSm6AE+hB4WkP4F2Xxt/a6dpUtPQmTlU
0+61KArBgOU3sLmsBtPTINY8cZl8vMzQOtMpHZsi4QxTItMiPXLVeFrGqauzJdHv
9bfspBt4vxYNPA26p+kEnKBWnNhHqvvG3j47WkSE7KZjUZHpFQrt5BrPWiDOkuGH
paF8o4vRzHvpcpDNgVT101/BGpUYGMAA0bR9SCEZy/um8hx8hLGKejCaeQ0VSTLa
UqHHIxJRupHhgqpNmMyTcIlo1+gm1mUlXlgGGo3ae1x1g1jKMKy0V4ntpg0koH5Y
Er8KRdlieB7PL2pCV/D4qrN90Ji06IVrh63ELS53QuHnWwXxyL7BODdiPtju0lKW
CBS3jN6r7Q++HvPVKFqF5u2Omy5BQZ2mM76b/4cxI3xLRFANGJ3zFWib1vMIGJcJ
Br7WT5SsIn1pAtTPEQSwZdJ1OqXXUJfak2pbzyrbRBWo5mjLs91r93CB52Ynz98i
ZOR99bxvBAuqFH64dWw8j5lRVvwODAs1HG+rPWxL3hPgkD5xTk1gO5ZC5A/pPpIh
w1FdGNJ+M6CaFUw8lX1lBpax2ZpRV/XTRatZMc5+tSxWPxySH/Vr0bsNEcmLFVWH
Z78FDLBXwkuvb0Z1LNS42rMU8r0CGTFkCdUWMAtOj/BdOmH0UQ/xWAKNGp3dcQNA
ifZWex4kdWXYhmXoPKgnJgMQtABtNlrW6AKm3FDvhjD0wWxkpmWQiquE21plPnV/
XIpC8WlxbLjpNkjXKkTTy2VauOebph+aLrlk8GuOQJygzOw65CSKFjS9aHHsgwWT
oH0yZC/PUdcDcJ1QFzmyz0nylPfa+mN7NxcSXuvZFTdcEtrIGdroXpT1gvgJPI6T
VCQKByT6oNEmGyu4Qer9+r5f/yZJXJ4xdyRibASa0YlXH5ic+pjCfpFR7EO+T2MV
gN7ISKnIV3nqMgfeangRYVdMa9/36I7QpYD7vUCu4pkDz6yzrgVjJOIuy7ATRScF
WGrQ5+zRxjsMWwMwWpkDhEtJixbPYgXmE8d4KaURF182VRY4sXax+81XlDXnkShS
sqSGc2xUdkic3kAOdwvPZCFuKt3lOQjNGCZ0Rh3nW8UILayy1wH91TKV+0vqo8mD
iA9qYmdkT+OXoKNFVnn7+D0ns3lTaXi+2hdJzqipUUT4ipwdOXs0fUD7IWZQZPdR
8B8WNF7RgpvHDWL+M2Gjr4w/H1OmZgeZ+ZeG/5op7baEQ4i6ZBADhTma59rpbC5b
pEKeehKvA42CG8J47ZIz3EVW+EZhE+RNRiJugOkcxiaZACWA6paHTCIuVlPKulIb
Lnx7KkT6YwEA7JW4tp0T9LNNlMDlcWRSaELeDfKBQfCasa/Yg36dwqbIS0HiN1Sk
z45MeAK+hSNmS5jNzi96inY3+gowcXjt7X+bC/UFpO/Sij7Fdlr7jWDCqZsonBfY
rRvCuhU6HTJIyF4uDQ2mKRo4DsqQC8ENocYDH1jW5RFhb99U/eB8jDhqtVdsMQPV
GdxvC2p3lVmP1sVj+SfHtNmXO5dsRw2Ig2FtqzsNSlYlGNVr0KQQJdu9scB343d4
JEMjEavQS9w68iLlAhvs9g00gGFvde2FTqevyVX9IR2qz/+fO5V53XkkAQa30BdA
uDCzYdArexed7gutMcLGnCOLd3HMb0gFgFYyT77c/6qiba1CCuwhx21tc5ukeLLM
bkLoFtyk5IBrYGJyWkIaOl64QX5YVVVQBLG3kTCkZ3QpJrVnBkmw7xvodBeE2M5s
teZRb6bxum5CyVGLdX5LXt2Ut6tWmSAi44cuCePIN1EEQ9kg1cn3IyRGK7FKanpb
UwoNjLtYO1IaTFohGruNswwKAAL8KV1pYoVxXLzxZlpxViErKXqbLVsRpttLxVw1
HjXGQlzhoIH4AxGoY0zLZsZaOHaJLPv6jt/O6jUY1OvuaefyysN6B1G0VPdra1WS
+sPiKgPohMSHJYsryvHazptOmufC1gtG1+gU/08bgXuIlNoyk46XXY7mmCPnDQX8
4g8s8ZjBeE+4+KdS5BM5ynPENVqVuMNUPp2O3TCNGyzuaJkC/AQ5E9tYKNo7TFdI
VSeq80xNCZqUolmwBCK8gDiZh2gUg3ZT1R3dR8qzm4ea1z7snKMxKpg4SEIVGS0K
0BzmYtBCvtUIE4x6YZMwdoKL5fS/KAdGdFWUfTYkhGXtEgz6kPmErhAWrk6VJpd8
38Tx5fT+y8JNjIHkdV7T/hC8RtzU6lqGewEgSEpw6xqrM4pI8WSPn3AYOyyLEmVx
tLlryt7/5m0XwEqgUjjMhJimF+rbDQueRxmE1QvnNNyaZ7c9Sjgo0OIFZULO4hXD
gm36xpxTvrSN+vW8cV8ArWQ2fekgogTc1CElY7npT/tBfSf0gad5JaB3geVfllEv
F3tvCedOq+iEOv54C4Yqx90/xZmmGEA9HgeOssI16mcUbyiZTLSW8Y5+KltSxG9U
Aou/UBN3CTtNbPm7VR6hJ3CcBD94O9kfjjI3Wc7tbC7O3F8Raj/adi2nL9VSoexZ
ACTq5TnS4rJFxu69Gx0qR6ysKZXoUnMsjsTZk9M9GoTSdQMXgybBZXuuuh5B19LJ
aZqFHNngi5ka+zCwA1pZesE51A8xG4cjkATGgCuwyHk5rhBM1cHoFPuRo+L1sRpD
FDRKVW6CziiRMmCaVQXpz+SaledJWK0xjOYDO9vJCMY/9owQnMQiZ9U6peMZGQdy
vSj/oMtiPdSdtZUezcJ5EAMgaiXVWfCX05cG8u7ijUsUL6heg8vyXRbJso4Awmvv
NvSJsXXhTMovl7bGpRpo7+WOAae8pITbVaACDWljJYHje6KkVZWnNYNd4HD570x8
8S4QMbj4h/pOjnc7Kphz8UNEOeoDVm0+AcBrrMzx5gDhrutlRco+2n8cMD6MY0ja
8KwaPB7ba/xrPqDkvUuEE/Qr4Cyw0QZvPSsskh5trEBwXOHoiGg5tjmlson0pA9E
9440DdlB6/qX7xMp4LTQhNpUD2vWWUqeEahu87GUNdVt+uNXBn/SUZK2wEbVG17P
/SSZusxg8oL32CHT7SGfppjIXzOPjSoPJdK5bu1CPCv6dwkvvOE3wAi9K2Y4wRUU
bcHV0naPGazoIHgYLvLx7z3YLSDodQbZgJeGpY/OE+FXflKcVkhrrS4UKQR6OLEC
NSzt8AcWn43jGaRlaPNDq8tm2M9sckBjE5kRcIwu7yqOpZHH1YaKaMyHYflfQkY+
M4HHLPmYrOZRldTUW42AVPl+lG2m9fdZbIO9hrzZfK/B0qib0ofK8UrFXyO7f6Gs
FmgF6EeRSoWvOziqsP6xojN6rC3bbyQqIS2ENQoezDKX/g+HpvPRgHYDUmpIvY4e
XJF4yO3Q4G2hL8UbIzdTFk0/MUG60wB7k4IKgWN90d3cQcsVMpB1WSTiZHlyx1/S
7z/8YId2dkMuaVtUudPGUClORVHvQ5saPz/6clYi0NrphcWxt5fwyjyI6b2w4HVK
n+f7Boe6/vpI7nyVsq8tgIrvTgx1eHjDzKeuvyAisxtkkUltnmyG4KgSoPbqj3xn
tiecqxSDtW7hP98N3FsreqG1WHLTgjDf2KnFK8OgsTxnu8WwhTnNR7f+XBEZiZTH
btidStJXvyHOKzl0xPTRGWPGbphBPn4OwdZvJEbIRg/XVnEH0fs2P/jvup8R4hgz
WfpMf9VmiXWIB0JbTugFc/QljD1FxR3btzy4Z5n4M9uBuSvxe8Q48GTKkOR9HZzE
7fU39cKYRDcxDCOptAn5CEDOpSSTmKCnamtW64auxnO2T7eEJ9phTYkHztZxL+dO
eP7PY1AW1rHJDJuywmOKFXtWvx4ku3O6xzuvh5a3MhVbjSjxpYmxfmsGzAVnrksg
3Caa4UZvagUJJdKO5VkgfTmQK2PxMo94o0nGJdvwYDcxFOZkbsHNFJ8d+EVi6nzc
aZb2RkHp53ZjGDZOw3otUgbM2Iybc7v9NxAYs0wfBlO3/mbgUCYzblJPXlw3qlmO
9t5qguU/ca+yyospjSxRLZTQ0SJDLXJlsZ9GHgjIJj6WQPBs1F/VU/PzNnk7kuVr
bpPQ9agIoO35NXbqJViIu6/lTgG0Fnb6EKsAMokL9zQm8q+48ATf42f2p5g7JQgw
Ga+bY1/YXnd7wWdAHgQpU/Ka0scyW527zmDmnRlHxPwDz9ZEPmOLPIqMnGnnPuRg
EbP4woet6I205Pd5MTtRpdGJOI2s7OcGvWSyInWxv1l/uwxo6FttXS7evlPLXtVO
fZ2NduICRH9LQanKUutFI/bNuD9yItzNc/Q68Pm99F0myPRYq9hymQtRaBsYIJu9
4FRMWxTq3REtCRORFrnpta6OKr2e7NCLcG4UMuKBGUkmdtTe28WtRPMPG7FpdvJP
HxTYPMCKQ0ErhtsZlw7sSSGKa3v56Iah7pmMmHQZkl6rDwPB6MqvdZAd78pgXiui
8mLj9chYn6LR1lcqrbMrrx4Yh2lQ0v01pmO2t+tDy0DKYb07u001cJynnJ7CjF2f
RyssODWlC6F2BWG9uwN8sNgAYqKIZ3DwySwD19hqit3FUPMkPEVYFLJKDRvt1FWV
ftUc4m6gD7IqTHNKET62VrBzAhZ3T5/mumRtMFtm3ZH5HJwSRpdlJ0ITmDRtKoze
Dj0aSJ+gEjWpV/AH8269RXM8YT+Whq0c2N3wpLO1AVrlm3TWRWm7GFfcdp/p2CAC
yYCb2tJQ1kf/2n7YaQdXK8mlxdacfJYjchWSLmrAbx+C9dFr8MqvJxLJRrIVtBq3
rO0U9/3thiUmz8LBsRT/oIYsgSn4NsjSDqQjfdZ7i+qJUqrG+uH/me2nkfp8Xyjt
vaktoxFwaGpXMZWlqtWekMUn9gn+tAFY2O2vewrriAdmdMCYIJyzhTj0lSiPwnnm
URQVIbJ+QOitnKgZQGEB6gfeBZ5NSO45Oz0Pufqb2oQISY11wywN4rVXqOpUI7cP
TB7zvhLB5BMOC4t3qzvlU6QWceXpVGAsDR3ODjuKsjTmO0AlHcTYmqfJvMW7iWMp
ChXFpyGZ+xe+O1KrWJRou0PEX8BI5RikjGxnYPlC7x7fbXNq34pwLbO5YRqxiJTF
jkwCmc03d2Cmup29IOh6HqzGhB/FxLpBUbLabHAtzdK6+Nwp4GKfJzWquLXnoiTi
W+CxZjT9KtwzpSDSvRqzw2fTeAwOMqAjp5DCw4jzyC5eS62sSKgBgnHqbI1ACk/B
cIqLVyeDjrw+7vtE8s6z1Nqyj4BEMBJ0VeCGlxpAhzMRkSbBubUUaCVrwQsGMGja
AsVSmIrcNToyZ/ocVnJ6kg6R4AE48v/s6fB70LdqTF6Z7WxjnFQ+8Tn5quW6wVIy
9VokwOA1uQ5jYE21m16mzoE4zliWPDpRPATFMlxub0JNcUUldBdUNqvL7EPX6W+8
WWdcb92WayBKTchbJ7xogPeuCXtW0h4Sx4KvhIoEHdXXnOYbS8kuNbm1P1NkoGVf
qTkzLhGM9VCKtEOzJmKds7/vJ8inO+GLVE5cUHVUU61/HEFaw21YXNGuJY/eFSw/
c+shZOOC88v9DTpPJ5EYeFFj98HqyleV9IbWDDFEAp37x/Qveh+/7WtBPtZup9fG
sqN4U2K/ZJdwAbR+FdIfmsd/0EjznrD/Ph3uWtNeV8EJS4HbgDHZvRj2xrYyRZ6z
/FzpM4pAoTkYHQ9gMPUF1DgPvTg8uOwPwhY4d0fouK5c7Eq+DPuhwTSFUwxkxdRC
yTCOHBsg/5PzuWOeT7nqoM8k2v64MBKfwGlCoVHgL7Xxbqwq0UOoFT5YXDLtTrOe
/JwITik1OYkyD3fN+Ng15Qd9Ljst6rhJKxZOfO/re75iZvczO7Bic1zXg+uCg9Jz
hVcyXNKk6j4QpCx/aS08Xc/NLG/LaCRPlF1iLvvMiUQEpNeCSRB3GA08uefvxRx9
ZHFfuRF+FIEzksry+n6mXqZKiXF8Zdl/rknv0fqD/eFzLg0ptkEsQaLEJgWGeE0f
lGYcVMxtO2OOQ0X82pYS/MPFrsJd5Q+MMbkhC2dR5AKG9kWgl+p5fi+Be6MGL+lV
0A2O2xAdbPKCHKYc7amwdBDwdzHYSuyBWUzS8GhXX40xBu/87ismxIR/0fnxl2Qh
++xl1sSoI2ujXuASPXv+CHWMKv9h4ROcLN8vgCz9WbtClh0oyEmYEttpLEWWGjDX
r6HOhevi2f/+8POQ8B2BCsXPNnbYpqwtdIAi/iuFY77091A8oh9b5QL0ulRu1gXI
JgUfrHmNVxRjoQnySsDn3ZJgssEk1I0zxk5EfZe3zrayh6Vl9LQ28fv9gp73YmfP
nTszeNjIeUE03g+Qd4hHIosDqyblEG8Bq/OJ08k1n101Mbt4yurAG4O8Px61rFXh
flVackSwkd7Gu/FECVubF1CcJ17+VOcHXWWp4cMRvC6Mke8JTktvmxOJx8HdND8E
n9uR3XI4xYJ2rHX/s2gj+isVX9eErfyV3jmuJrkDNAjJ0575I/P4bk2Fd0tB10ja
aL30pJfgANepqD86/pspZmZzoY1idRajVUGitZeM6Xa27I+BV0ZbzpxGGBv4gq8A
EhfuNGrekYU/W+mJfGmi70viCI7Qc7SSv3Eem8XuC8wZYqXOir1c8eq4opsMbHR4
jJePsgfYtY7D3y86gMfOvsHjkdqsYxFMSJtAMMcJ2s4x+yLMqmgMyomFBrOAcoat
BFC4taMFWvDUQImL9+ET6VSNwF3HOPbl22dVx6AXMFigScpMJQq+yfLYBagkliGz
iU2x8b3u3HmDNi5DStQS9WHFTcUxopcDaIIeUoZfkFrJhakhyi1OHEfq83a9CHch
DHKrm95Lb0qsFqfRHpsW066KUYsyeviLRSJwYFZOfwcJe6rEEN/32lCNQc5ByjdJ
4V17r9rlVNPcvYPqiUMTo+BNF3loy6/4/z9gN5EUAoiFaUfgjmkFXPVd7bnqv2+E
jLXmIM8A0xOzQoG3RAuaXIb8w/mkWClD/HAwAYdbl0gKxKeeZuWN0UqQb/nezsPu
dyGbdWcxZxiC4XK8x3QA3p4zivfWOjbBWEf8cp+mL7HINWjJAzSsalpfQEBRphkX
dIZAThCuoCWOOpll11NKjwgxt/DeTw9OA0Kx9pjaiW205qJMMffEh70D1DXIDnJ+
zZG7xE/Ku1vR8qxcxm1ryOcIRVeKpSmY32EzbnvK9ftB94LhzrWc9xS1JQI3ah9D
KNcNJczmPVu17alVxhzZJxCahZmOcQBIGL3i+cr0T0m005L89JF34GDdKj85We+8
/RFStk16QKHQDAKhgeEItXlaH6+W/r/yWy6euqPwBiYNPvtqOI58fhy5REfUFvpG
2wJEPcRa/ujg1QjK7HWjGRP1swxjGAO1eEcMvLyQYDXQrZeRe5OCZZQbXJUa06fH
zlmvAxt0iFnBn5/kagz2n+O+xEAG8t5jcnrFqNt1bpB//A6d5o3bvmcbB8U2p6u6
1O4dJj4EBFzABpEq/O6eQXdUNu4E/Y92v865RRZlKY13B5jbYJcyFbeIP9KhWEi0
BnDwuxT5MLBKREBRaBT3beps2p+3DxrwwHg6ENpzB22M4/9UL9jq9SsBoiqCpYyp
RsnHivS7IVYY/JZvLu39o1MnbhIADkg4YF47Y9Fh9Bzj7aZDdRwzyp5Do2Cm2hEq
Gv8WuIwU9pice6xg14RvTfS75JaC6yX9BnDFJECHee12nx/aYw8KQJOdbZKKmMh1
FS+G4sJx1QDPlvN/pNU09EVGggZcXmeT/YrZ3Im6/FuIKPm2fjd1QCwK+o/hxZIu
cyIbGSofStpqTEJgxHq4dpJVMMC5cwLJI341TwM22sQM/mPH+MhZ3ZNBuTgoPIB3
FYTzkNdDTzYlO03hKvpeuG7Ry9U20A8aGk+Dxn77rVTAkd/Q7lpjPc2OeW8D0PHX
uNNsmJlTw6LXxia8BFIUZiPrM2HZCK+1pB2VqfzG7fYXpGaZqH+DN9Gg0fpNoCna
nWodnR/u0SE0W7VYXoMz4cB32KNBfDOhQQC4gIq30pDN0vKbcnQ6IjA3TQUbHTFH
XnvPmngcdbzHNWPFMYyg0XrHHxkZIIwzFynUuzrh9oFD/DYyPSZe6GJaWu7l6lUP
Q2il5QwW8F1lFjUG0za9/Ow6cX9rAFBmUE9faTOrpa0oZ32VK383DkipcG9RY/7P
F8e7k2XkaSrCmAvtKMvUwF/q+dpG1T90rtpw6FmCg2GYvZ3810VC/Ffpv3SxQDC6
LZ4FiUaMIs40x8iM388Y/LEuEKV9V6bKx2lesQeqIkT2NdxMRmx0/oVUBLCyPkmV
vc8Y12/a4i/5BaNlEp0EaGWxaU0lqPttmQ9kOD3RTRiBiFX7DBscWdjkaK4P3aSh
XQ0JKuyWLtR2n36ytE6bWuMHdwgAlTm6J1YSAenNIPXBdafavluhxW0RTro9m1Re
8HkitfCeWJjGSaXrTDN2MjMjbxFyShKLohYd6OQXxcMja+sMBzdThKy1rMSPJC0H
vHrhZWnzFE3QlbivrQ2N4I8enqak/SeI65NaIz8SoeJK7m0mEN14pmvSz7L6hc34
9MMOeO0YcDI7NAhcnSokxmXZ09kXmRettLZQtZFwq189Tlbst+nQbAvjLxfGXmVd
qtFVdvq/ocfh6hWtbETg/Gsv+9fOaNkueawu+JkcTcLb4jeDfDWvyjC5U2XhdDtg
hqTD1bu0jIf5J95+6Vs3NqD9PD9fsFeJLM6MVJ4OZCPX7mXDEEvsvFtAD7pz31Kl
FQ4oJjaRj7QW+/ThIS1nbt2KYY+7hj4cMSbEqE28YuylbjLii05aS5fbkXShmfwd
T/BV45Xx9Yi0X7HrxAUdwDsMaSVswLoWFl4nQmBmQpdpMc8pGaso9HvezNnxwo4P
AWIYphsfJ+WaYYbbSe+RLicfHYY3sD6wN5tYYnzyeREwjZ/BF8Mfjuco3lPIZukh
hjSWW+jjCNH9WyPives3ZlU7EdpyU3n6wE+qTwvCxOtMXlKgDMYWDNuc9SqXyIOy
iVXZ41nQr8CrbCu+2t48MmbbT6/WSBmYlToBGlVemjlJO2uo5L8u5SK6gvp11dmU
ODp3sDTLSgeb6oev9hSqEWL08sitIIYuCOfnV/dWIr7Cjcsw/13UiE1dIBdSw785
uk6tQgf+vJVMFubePZBvrUpx8/UUnlcw2DKBHb6a4WJt7OMzm0z0Qai8s5B6maXp
mBHQqHtpTR2Vue4v2nBbPBa0ehawwmZFhXoV/jyrgC35M8gGagepcQhRSNS7/6XS
dn4licBL6F7fzx8OyHVVT99CcqSdVBNJ/jrUfqe/TxdR1ZA8+8K3FI64/BYo6JFB
KeQ50Avyk0Vkm/30weD8LTO2VfV/1VuCDg5BBeWbyY/VlJn2vhG+VF+WZYzwx5uY
dF+rDXfffoZ4d1oaR1N2WbOpapyrF7gdQj6efxhU3un4QA7qNX+QDyR0ChYw02Oh
jSAcT0UvO+r8kqDB+ZJuqu5Y8m/SNlQjbIJbrqQYQ8C+Or8OLTCKt0a8I0Z3FIUC
t0BMITCqRv54rwzvDaLRdJ00fOBGt2MAasqaIh0HYS0wsxsPpc6/HLmLxCXuxlnT
wqhsZ3Pwf9i9YezHS7KAcv4GnzEcw7KTNgU/n8C9chZEOHY16BLwDx2dXcARgqd/
N8GlnDoDzAYR7Ou4wvoifi++SBbjUnidteQ8psWf+KZPnPH7Gs5l0qYpddeQxQ0c
2eVmn2L4f2OlPRLe/fLsrdlToQBpPUmPwwXAigveRtYbNXbh8W2dc33q5gRmbHow
UrpOEMz4IZdXKSOMiV9wfcvMzIHIF3rVZXIFJ0OW9bN27iYgK6nDg87a4MwSjWe2
TBqu9uZIirhAz90uuE6/ESRtwFT1BNnvwjk4QFal/9oNowiNuyk9Y1lSmWchpcky
hMlMuwN5m5Oz1DWyXXld4nLG8YR4jCJyUjjkla3vVJJUK2h2GPm9WdctyGbB0myj
UlvUaR8AMCCAdZw+by4VW3fpZpRe9Ca2I1rZYYmW4wRfWa2OeVzkiFXpZBi0rlMe
uxe48hXkVFQTcApw+Yp1O8oYT2uI4xInqwG2NNS3dHQXaMHnPQ9R4wfQA3nkwO9e
HqHzX4dO30bqvTMWXmOKNfa+2xiNvGGiCqgW8/U0EiWjY94RWGe9I7H7Th2RzZlH
GoltcHUGJ/318VRIzgNzSx8FWRJ//V3Zxlgckp6Z5Kpb7lSZnZTbpKl7281utUZb
rY1P8W6/NJ7BAegHIQjFXiryiGOFqXyTNzM21Nhr7Ynjy2vQH7cpkeo3zJ1LudyG
FBldgwyHGxLs8nlsoZvq/yiYQabRl0tuqY8rrjQZ6UqB8p3YVInGE5ELdDF2Tjyr
FKq2hlHyicPJ01uyVnaeZzCcur8daonlWFYiMt+lj86zM0Fxfk7a1WB3wsbDRJ5m
eTo9EPgqMuJUgPIBsEJOS2RHAmMaob0xlKw43wgseqHf18Tibrnyo5NJwklmvKOz
bo0Xb1rFhivVw2EQwiZRnjEjsksyfS26WU6XRIEH14BgPXeVau8DXrwE24a7QYB8
0ppPeTh8egMgFcGr+0t1y2dzvh2j5vpzMexLe7lSZraG8PHYuU1Lx17bR7PS4ZsB
gjeB+FoaiQY0Fvjoza9lzByAc26oZXG7+RAGdCEg828eJD1LZYj9bFyFJp2onfNQ
q0g1/uA0FoLrfQaABmowSyTJK+muGTy53NRdqeOpsgYMwUyDyGiGcHY3fyBnyXA5
O0KPXzjv2LdOArZoYe29s8we6AL/9hhXhAcPLDtlMBXN9hHmusQkbKaptBJbQEeF
Ixt4GS0HHcRiiuB2yV6bV3VDic1CZctWuQ0mZgDfSfEaN8WAg6yD/OiL+y3rHaxh
Cl7ASGzBGpgW/QxOCi4QuwGSWBoSBLtRDD8/+gJLtk/vePrD+4pZ0Un+TDQe95dE
GHVzDdK8st7PNuj+Kfmme7Jvq4xzMvzK3pYLV48tobSGdB4OEHG16L0DhvcrnoFT
hOXr+u7Ou35UNuQKfLl53vYkXRdWzzk+O3WWV0LqP4JpIl5GyYudTXSTJKM6LtBh
ExsFTCArOBmrISrKU+s6mmyT1Fi/wiU8vl6Bjk3lQ+oZP95qrhRnEmlVngpEv5qI
BSF9DddbrDtA0OvGps90rhNUs1kktL5m9S3Rzeq1izigXEVNjUBeLJ1MwPAv2FXk
+ak8c6vnGr/WOTMm0S9XN/QX+DNK85IRzAsPqjXJbYlpbqyFOBiBUBA704Jf4e9v
1ObN8CDT568efLyuLG9bRNfnA2p1iN605FM63fbe6XgsK2CBm4qwjDkZml+wJDAA
URk6LH6AyYNwABT7MsyObWNxxJE2oUIHtYtjGIZbJR2Wh8ZsbSImNddKKU2hXkNE
WRprDpX+iPdmuDgvh48fktfhkmP0Liro5K0dPW+HxAKdvBkDK6VhR0di1VdJcgKp
zWyjHCRaBs+QrRYaBtMHgs0ez+kwGGum2ii7kvrVFt2kja8IlJgGWZOA/IAuBUAX
G+owRHMCDGS0o7ZnMeqTclHfDm6flWtekJcFDoOLDVfO2/ylOKXhU26GjTSpioi9
OPE/OdA2H+ZAyuuMactCfj5AzPih+Ni6Mff0VGLt5PkQRrvOGDonn2N4lm+3CCN0
7zLDUn+xZmUMpkEJ1olonB7AZOEcRS/OR/GluUSO0h4P2n16byfdqG9jyO6isKHo
W7JOx5BsGQaAid0g0XQS/kZRjI/Lm+VGOv9Cgq5TxHRdFRdeQZEpKoBE7p1fkl8L
2o003Zu6xL/rvn59INWynxu7gzvL1fTcqNVS6S2Vgxcc5TXnuG59htP6DV+1V0sm
6HVfkazepdSw2INB1g9WSxOzcj3nfkybLf3xLLG9czpJvQkZMTEl+s5s/hLS/UbB
KRp8ecUjeKYNDf/94eahaI0dOIFsaO+Dnd1DTzuxQLw2lcWsm0/rl+nHlBMoapyS
EwRhmD7sqx1LoUCw3l3sf+LoFS60SKfh/aoeHdg17Pgbuzo5RB5hiwzq3wPLmHaX
DWwVrUwJXirTubjnkFLwohhDJRixcpAYgVPnSs1K/0SmOOTrgGp7S9qtcW05jZJj
4PlUjTtl0qUkC6Jx+5mfMtjFclETFac7/sECWpx9XiVSa+QOAzZIrXHbmS6oLaGQ
WPEr4ATN19g2dtXmpDBzhrROEHIBFcij/WzRUmBL8BynPpPPGY+ekqIQBle1U8fR
neb+yL5MuniazcCrv88vtFFZp/tuXsqHKCI0HZypwgZY1pEbqm+ZxmgOLzJM0GkD
e9KQDPH+KAkpWDIHzuO7SPJVpA9pRJzP8HDfLkjmO6EoJHzLLRukj7z7nDRYBG9j
98f2JCNHdamIM+M7NLPrAIkT9yTM7itR6Tzf5/fk1nVYK92fcHz24tt7vAyAIdjZ
s6vaGReqw+1uq7nsxlGDH8npDixZSfynCRv+7rWpBX3HI2T64UP0cmQ++iyP1xpH
jfPQnJiShiwUbsmjFWs10CrtKew4Vg18lgTW5C8NZ2sh0cwx4huJWIxi2YaciJp5
eBK4i0aP1auMh7I0USGlRVaJ2q1kaWbiwGEZRtdAN+V5fKQdLLq/xQVO2ntiDbyX
fwR9Bjq6xUjOZ+7QuNfaS51yQ4AZzo3vkd6T1Qo1YjFCLzVWQwX8d7pfKbghRw8b
OF+ZuosuW+cNJrSQQdoORU3iTQkG9Li2gzb8D7NE2x6y2pFRJObYf/e+BFc0Ilcx
DNYhQEOoGQ+y/yjpaCAxacpAYxEsDGXA0A3uBWAlmg55zFAa1U7t0GuRYA8KdxEg
6CDN2u72M37h+W/bJGjrTtOwLcylDV2At8xh6zApdemaIka+pJA/Lzcjhay/fp0G
1saG5G1KqR8EAFNJjf27u/JlLxXUBHyLEdYkgStWR9TlJs9v6OE4iHwU6iNOwxJ1
vlg3FkA/KgD30a99xr7O79LabPyj8leRhd1VDTCYsiwRSzmQsbGXTblcYgn5Qt6W
4YD7GS6BXJGm0xfnUl+cN6m0IwYYCvpb88PrB0d1jW1HURqV2Zv0+NLt6/driVQD
vgIRevFdx9mZyLGRMBuNOi1jT+y9oKq5QGVy0vyV7DPKSuq2Em+K1+iXaXXyT8Bn
5OQvJZwBUpbwFIZMl96e0xsueICNQnL5tShSORJBmX17eN9Ytdpsat955ZT8iInB
DML0FsfXghAO1mVaAVJzgpNKQYnHWSU2H7LMwTm6WjVXKq1qtqcB7RHGGSwOw5Xx
bcl3lKeaXh2cIw/tSA4FgyVUL2zsWtL1cJoEroT0qDrXoCEWo92LqX++PaU7y0Sp
QIRrvBoTg2jvv0uNX8onvGgPjEmNN2TN8v/hYn4RYcDA25nDPv1duWaFfbUuHlPd
ShwMI4CYi+XBZX40vNdA8y6EmiC5ZWBXI7Hlrd1enyB+dy0yvYEsqRR1CDgI3OZk
Xz7ypnnxRI50/bfvnqgjcwAyl2mIMNyfk195/G1xUAKcO9K3ITskGQQSrqIj7W8I
ejIJnli/+oq9rXcfwwvAdrzFnHTxGi1Gze86uB9mXlcuap6AkkoZkiZ2Srp8Cd4z
4Ti6/7ZGJlA7tC8yVTdy9xYH8NGMcKiiILRN3jmm09Zi0h/lJCaOAu7UBUDwvFGw
hLVi6AepFq2oa2+gYUqtjf0ZI2Im7nAH8cPf2Eru4vSNjQa5YofrgEhO7BA92T8g
togF5IqkAAim/M1NiCYLdlp4HPDI6birEpo6s1oRtASD15o5sYy2d11n4nOobXTR
DQYT4mvkkp+AOC5dU/iWTT/6KlhDT6f/8LsY5n+Kduz3DKOR3mRDrC2cvje+MvVi
P/SmlcC9LucQB5Nok8rJ4kfKIKBcrkasFgZwScwvruDoD5sT5GFMP98EX4JAyZTC
LBKLYO5fLItwHbRYYjlji/++rrgRmN8CioTq3YIFXhtAP1utwyGlylnm/Ix8/6Qd
qRKA/pILCuIyxN0N3Eo55/xD6WTIp/2SZ9tlxwoGdpIXNCH4FQlj+NBzw1kPxy7v
0f7veFL5mT2lr4Bs++Sp7+Nc8vL5xLoi0IMUgQcJWY9bvmCUDghhXdjdTY1ufEx1
CmwQbRzT2QlLT/F42PW8WtJx64I3LcEj9vpRU22VPGVlaQ5BWRStbxOkD594YH7r
od2II8gN7h6uH1tUtmQwo6PKK7RotIokREn9UuO6nwO8zQ8EwPyOosW1stRfgE5k
nHun1/nmnB/gXbCAb46KLgxNHn1V2+wbLHLmfxXvVHVrYjAjkPyfSs99dwfavCMY
6RA9DYfImwmMCsb4D6i+PQCcpPJGPYeuWXfOCaPL5m5m1DuZn36Fe1lYpfoQQB3k
7lgqDKNzHVWS7VbSa8c3PNwu4RxEVt8OEcuLE0O8B87rpKriL45iYz/YYuuji3/G
PE4aqGnsunfcYOV8rDIn2V3ySfLb1244/crY3DCqSm4C5IwmynfvzjyBBpCMxjWw
dLQdGYJSS5VnCFqfov8znEQxFUZETmzBaJBiyrp3D32Q4J9XZfulAA37Tmuh7CaN
6aiShiTBtj4shIz4Rnk2daX1vCnduJxs1U3Fv8XJjoaqZ6YTh6Di7PUS4PGgbeVv
GfyQenpHRZRE94W2JN/ydR0T1ZlePbZNg43k5HqbRB8knLttujS1esf8/koM4BWs
ZDn0//OG64RqybOsO7vFqXrB2CUmOQq+72vi1PgFNIzqsJPriIBZzsbnokqnOInd
mvo+TRSVVOOm8V4n7BNJD/sPlHPbnZVY06OtquF+yzFp899D6/16Xpc9n+hlE/VP
he3M33d82xV3bXZcqyrMXb9uLNu7AUaxA8DZOiBRaaBrbOkl9foxSGonbjPpuPsy
wdT71GMsIciiNzyJpqE4pkl85/12mS/n9SaJ7AsH1k6NN7MF6EuyVmqnQEoa1zxT
59PrOa/yETy5dOgsMVvffUqlfMFQsl4GgbnYqiP3txpPGKxNnqVVbDDAwaK4JpIN
qmeauxN1Xz4ECrqB+WCvVmKSB9oAd9Xwj6BaPlY9Zep2Lw+6mPzWr4qiz8a5Zi3m
xsdY/fDJ5BLQVW5rr4Mrbzr7mSZ1/zQAKZ7rbuJngeoZ/nnD9rNhCcdLAkFfSAgI
aIJbEhz4A5IBm98toJ3lIl+oT9zZ0hEoCqXZGg10AnwSSMqweUB1zti7gZF9xMp4
m+JsGUAo4KFbluADoo72Gdx+6KEBpB5wtYbLLVlIf2GGp++J8L2EYQrKwH9DVgyq
73LH6pHPiAiGfrPXNruKD/f81uCR3W1VCUlHfg8rBiqF2m8zmORwLn86y/vqDOkA
mBHNU2tuV4bWqDP/TAVfPb/xocGucHemZExpl1V4b8mRDirpKiWwhl7U+LiQ0p7A
QquOieNs+voMDw47Fnsgmi9fr4coFhnPv3/uKyp61xZJdQn0IHsul2xAEYOtXGhe
siVb221dvGO5p4GdcEHDhFjNncY1r4zzTggsQw42J+VyFLX4NF1gzvKMWgDqxSuA
LOdu2iTvp7PMW/PRW2QewDzqGgQF40YpsCRGQBrxWtPa8wkkKKyvZBc96svlMmSG
yW+nN8WrJnZ8iarWX3l76n0fBGJC8NYfyazw5OjGXDf1XTff1bt4lnUwIkpHjLbn
T2D3nt7RsS2+3HI89+J+xDIXM0KDiFVdgafUfGZiuuvjjCaXnqjChuJ9+rK56XcY
mJPoUhroZD9PgerTvLLXpioODaAnDiZ6lZpW7t9aJBZ1FpVBe+B3J54KIet2uyK5
Tj7qHem3TORhsdM62IhYJJ+loQv5AlXXdLbOFgLpZ3M5ISdpYG+UhYH3n2gjZI9H
tpLYaz1LIHjyT2hliyzFOriFkf/+Ka+tQTz15ajphtz7tbqt0OC7H4JRcLrIxxVI
KFkZ5ilTH/YPwXmv2BqnfqlK7/Ji2HFPuRwT0VE7f61vu1WsJ2VIEuv2WLAZe3VI
cYKT/QpguddMM4MTsU86HRELrCgbAa1HgA5sHPsvmQQUA8qgKyX+ieKfglenjoSN
rbwbsAS2sETOa/CaTzDK3a3f79Lo8sYxE21gaXMe4XqRWkWGw/BLaxTt+MUX2btH
oAsAJ1zMmRPeznMJBthdgX4lnu7nHfAJHDQ2DXsnTTeA/OIbcMHUOmGH+wPSDw91
O8qlUJUEEgTSLKCQWu3Gr9dMQZTKPStmNag5qLfOS0IL81vz9lJWlPe1jrzZF9lR
DlJOVmST4mY4rEXe4blk9L45jGcb6KtGsH/ZcxbK4ZsDKRAoJZQSt+xjTVJ58k57
I/+gOX41DuxLU7uCB86AZrj9Solkdq9a9/57UkgY/oXzVEgfMs/YjMWC99bcLUQy
X5DIRHLHovrrcMs7T26syFxZbOWi5CQ0zNfjhvJ9Nd8q2SmjWt7066msjZ0jVSd/
W8KH/8muU/+zeHdDRC4lorLO/+HuLjCgxOENfs9CJg6q6vX8Z7CqDvpTBbQAbYWH
4MQBaPMWcYVDB2Uq8ALZRs+mbHwdY/C+3ckRcPw5uxnUn3Ua/eg3nDj3flWbywUB
byuhCgGe/rkL0lMyO1xpgP+6XCUVB10oOMi805Ny5A8LqmsDEbiSJiwNjmX3NZC+
BNUUHnJn2P3kKZKazWNEC2Bv6AxxTesebSMroiW4E5D1EZ3Urzx2CD6VdnMfLjnP
x0lsFpFP15129vIsQnV+s5lhc0sNKbo3zFaJ8whP5ybBssjTfvQbaus6cwfpWnT7
UNTea8VSd2q4lV7t1b2WUhMjYon4AYgKSkK8GTpSsRn5Jxse5hvzcQGGJXE2Cz4K
ZFW4FKDOwiMLrCyg/w1wTkB3v0LaTW9KnjyYhI3aNTSFlXCFgOV60V/oA5xw4m0k
njg4firCaQjz3alOcMqreQNOPBoBbOpgvY1AXlRaDRJMPVOAtSRapblkdeCIl/To
UI1SPre7MGZ9FvEtQEthQGffHRd6HuGfiO+uKgfo+mDbmSGluwC6sA9Q87xYEMyC
Ypsm0d7HyAa7XoNm5Nmfw+UBfvyO2L/o/zMJdM6SiLZ9sk7t0K5RnFyplp1LCm7q
XhE5ifvwGvzkK2m3OkJU2cNowWO8xTmDTL/pG7VFRS8Egdl6dorLFdG/FxQCzth1
IdbJIy3REQMGNeyyNjaSe/DFfp1oE9a2lFQyAE7Zjx4h2BJ0WXv9RRK39KuQFYnL
HmmRGsCXnAdAaagYrCh+BivAMFvofALF2MEQosAaKuXam8jdvU+RpK1CzXYJgvLt
ov3MyyYoRUZrwhcuYx2+61QH3fCChEmOezmVHQDJUWoe69zQ9scfRxX1VDJ9SAhA
YyD9PvzHM0T0WpRkTHO9dVrCDmiiIK2wx8xNORoLHmsIIv1REm+bXVDya5MHYSTj
3/adKGnbn67+2uHd+vvMlcaEsiCYjmiRmMeBAAd3gnUyZyZjwrg8Az7e4mH7IZoE
OnRa4wXRnsZtRA1KRODtRUDZMxRysv9n1CK3qDaSt2pTjcPqWauEZkNg9/vjtcwj
EQ1eg6nHzEXZP3MC8zCSqbtXwv9f0YUOR0GpPCxADZSwgeEGvBtf6agQoDbasX0T
PoeSwj1ptz5Djlt4GZj8Yb7TyfkMm7sKeu4No2Ezw+Ye9MzMpmFIiOVmngKKzX80
KPWZ80zlwgrCKCT/Pn4DZjlWSxW4KLs/udHLIprKOB+Bix7y8/W0oYaL7MgoeGEk
RPR1SfyRKjqZFud0OuWkcQcthEpF0WRLJJLoB4LcDekSSiXo4PI9Ysj96KpNBryd
hMocl1s1XcJHnBKugapEDFgpuP6zKec7tKm2OE0fa1hWNCWvT/WymvfjmQqqTzB0
CbebY5/SNtJ4vh2VZePapmjX3rFMghvVwfZAlQ2XrNpQJm73mi2kPHhHgEXw0Bne
rAYsZ7ndh3RWnT4MEzVbHyJyFz0h5xpOe+s6CbvdTD7PK/yTwX87HKGM9eZdHGsP
R6rk44UgYHdCTb1T7jvu1xX/oIryuWYtLxAEeeQ3D8o+nNxhkX6D/ZtfOn+pj4kj
V649MHk4yYc4dxrHkj17R4b9CvYhuWRNA3oXzxcYQluGYp8daG9Q+jXClWgJOcRB
fuCOYJwu4sJMMeEO/AGj47zFDv5rh0ihplWbNbh0TJSn9IW0ciBzfgxDnbM6DKgw
0vhNULpAUxQhd/LlWyXBuBf3U/ISiLIh1EAccePoRhtzbjTtd5JYPQi67so07dmK
t4vYO6SPLPiNWb0Nau2r5kbXJakpaj+TOp9i5OcxbzFcoCcTyBBuJ1baaJ9VMFNK
A9IUQ6kGxSQLw0Q3MDKHRWEDU6TU5m8yDv8bBgoWDAzYvnui7kQFkVOYvYAjSsae
NMJvYkUlhNUr+J216FTrM1qBgrtBfnQ417ksP+7BEPmB6Zww5HnzmSCq7LRtEik8
j8I0YcldvPwjixbAnUGK8hwAgzMoKl7lPb9Ofj2TlNKYEypY8wW0LyOnMTmVZn0N
te7LA7KfASxOM2vf7QK044+YT56Q/IpejASpY707ivrcN8m2apccKNG7yp/QrSi1
XM0NIGC4M87cnRiDhNWg8pIdNmmA6CgF6xgtQhMjP05zzS9tfibzY+U66WLT1fH/
L8gdefBhxrhbldVeddjwsgEd0q59oR8M/OOE+T2JSOE5R5SpcgZKzwmVgM83JbIs
uppyOn36y0xt3q/AIizXV4FMI5uUjFv2wXgBnbQpRbP6/iR2i3P8LBowrgZ+Df2A
Y7UnQCW38SUR0U/DyG3CCAFyJDWpDd84G24R0Z9XIAuWKwCjRmBsurXeDuYzTYBh
65qkvK5nI2kduL1vmrOr+S2Ox6s1/oj/Ti84zs1dWTipClET2oJy56hVs2kqCNws
JjUWqaCm06Jlvjk3DHp7oWt8Bcsv+64+B4/oX2ImueYlB4N3kWw1rs0ol37qRL5J
xJSrJxxkiIIKxn7zUpkk7CCTwotHzpfZlhxxs5I7NuR4rtUYjXnwTKvzZ6dNxa+s
0fRZGfBrA3+Z3L8KTOrxYBdBE5qva5miDQVBTTrOcSDfQMgzbNhkZP7SmSaLed8t
Slz2nrgZtDpVhe3msIY+jleIcSysLCNvktB92PHx2cOWLgbVfJFfRSnpPtVDRcOo
jnpgI10dBWx6XruUv1qPE7gZkBWxoIxhhB80+qEmhE/Hfr3UhCPs3RQvT1ghZvTI
6MQZrA4cQ6Cs12dgEebBE1Kj3Wz2IaW7vS3QqKS87FANBV66x5P2+nO5a22t94+0
JfOUAIhzH7KJM+RJX2f6dhh21Hkkp0shQnTAxZ9fXbOkE2FmYhB6sX1cz79G+oAT
+FeiJqICD1YltcMO3R4+AxEoclLIr+XUCO2dFMHeYIZ6sQGarq3fxT56/Y/ZGnhy
nTCNvawJIxMDoaB2nUUCUoEi+MfbzriHW8v8uvP+EJo9GBFwRohlAN/+JZRStV9l
6j/BZqMjlAfo2CeRo3ANKhZeA4CrEg3t9aY7jNwbXkx9yzaxcJv3U4nGpcxh/vyQ
cOMoxVWocCbt+eFLCx9gpiFXzhvme7D+zaDSz0ZPez+I/pMuI9g8/BvSCL6KjVcU
NhZjnUK4LYDr6sJtfJOfZD8vNyhGFHt5mb4T19fxW7VZ/1jBRXjiw8ylB1JATAfK
ZXAVjeGgjAvWM9EQeAKso00B3RLUJYdv89y+0rOE15xzrUIy8ygv8aPMJiyGAhcZ
rBDcog1wz5TqlbuJNoYtvKgq1OyoQZIQaAmY66zkm/h9gWTuCp0Re845WfGvM0rd
O9LvD6gN9ok0RpJWjsIQ64S+C8hv5Fav2JJI6xxLlgnXV70jiL2duLMie0hhCzir
xl8TSzQIV5sSAnp+5bKlVxjT+BU8yIGFjBucJCRUtx1M1L4RaIT8yskbpYNi6WYT
0rHLjxXGC65kNfdZtuSmh64clzV+FMD34oYhh3G7KIc2ZNCL/x+L7JEkgwBoKN9x
54ITTGwg0U0MLOMh0jG5dpJouOt/fCpCXPIYLJqiL7B6ydK1xbB8HOz+TeLaJOgr
LjTINhitRwxK+OH1QGamAf1pNfaruJDAVgf0yjCLlh3pwuFPVhfsA20A67aR0gzr
EsLx4XPHOa8qg7JqMBjmGDCxUk3OTqnR9bggNF8bmLdC6bilHwZRar8tEVs29bfD
N3atjhZE7JwzgciLdFBEf9CelMfakoaMutXFDSng+vABfnfCsOX6+5y/PDpIGnJu
J9Dwn7W6q6QcCmafTSmseVPzQqF9Dxj7Q4roQ+D4+Q2EZWI1rPbwt9BbfskBZnSP
PyvSWo4iRmZqacqGjICFcOx4N60UnQm+NeByFef2oVSnKQTOE24PVqtwXlKD6PXV
2iuQ1yia901z/2gmobOfBiaAamC4OTPWNjjqN3Y3r4WGGaBwTt5dSw/Zm2AACT2l
6mn3l+KoDkQXuuPD+dRzteTliq+fpd3KQPf2WU2pphgQmh/HeWBwvx7DozSSwS28
6G8lJWhEv/erviDvO1rPY412YUko4c3wd7+F/fNL4HkcG3W+45y3NTvYJfWPskzf
7SlY5hSiL5jgX+dSAnVazmYvrgr8niW9theIq0NbIEaO+/u0SkWzDCwVA+L5xkCo
44g0cvJYwCSGV0l3ejPCAzajvjdAMPF13WFR0xGdzwrF5Pyf1xeT1qsW4tmZp8Xz
aTyK8VNphZf2LpXlnBtpkQM/fGnZz7RzGjsROc8aLE+kgYgA1K4jvAcEoL2VaG9f
xJFxNXwifXgxNqYa39Qc2fppBxFUgpnOGIVEi1uH/QfDPHRxT6yOMuKbv4VCfhP8
rmSv7AxRMlAOUW4QnjiwSbtc7xvfWxN/POQXRaLP5q2EPpzsUho2Zp4BDaDgZbOv
MOIg81LP21r8M6nM2W7iM2uKmdwuP/Sn//VTRTNGaBe0xgufbtfYvHBq6ilEaeGw
W5VM8kbT8xcAyaO5Y4r602gDNs0aZ/UbgUs7du2A7GLmsrvdrg/BCdfDrp10Aak4
b2QkDXZxiKFb4nQFN+jt37dtsFbajW0orQZkPtUyWpH595pQnfVKVDRywfc6HKQz
9MugePVZ3hx1chVlaSgLitgvUEca6EO5Mg2JLaT+JoYTDb3zUCnOTd8PvFdIbzOG
3Jw1nsJD+k+fd7XyRljXNxd2oVYb4FFMMxmuhvtnN5bp43DiGRvklblJbhWiUEgB
i3ox4tXzmFGjwfmCfauzSeyt8rdaHisDxCgQG7lMDXYcfodIsl2/4N0/BlVXijTZ
mgbMbhmpvfBJyXgfNl/gDXy85E3LQrhLS4DVHkhUQ+q1f09dq7pu+cQMen0qiw/m
5fQpFbUuMODFegGeBhHWH2aG8LtyCyod0OqBJ1Cy1VOFkwi0JYh+RavuaBt9bqLe
48g4MICOHRPijf8X0ydSoX5IRr/ADOpp2SxZEBkhIP5msENqf9XYI2TmQIjZ24Ej
rMSpb1wn0MhnKcxROlZdDha6Ej+/p65YnYWb/54jDlSJ23T5EjqgGvFwvdZfW/QQ
NIaVontQQCzEuYZCWeqbzSe/x8OEjELGbKJDa3W21yaOm6Vu9BixTRfmLoQaNMFt
jei2K3YKYzhXc0PB4JbjbnubNr045dp5vnr9E1/dsB5HywT//XaKsBzKc5LuAo1k
tgQdf7H2ffV6KN+mFr4oLMYikUU8TtXyzdt+FTTyIeLb4ahvQUggEnNhDLR1bCX7
oQw3gZF5ZkLG/KZdt/lLChJI65kexdvrdyqP7QjnuWTanf8aBBtnc+ek1ghJufrw
LzZnZ9VcfkCpPWYfPTQOryOCFMHterRZedbHeNhDJHeK3U+HiecftHxq6grJWn7x
7PGIX51jnVMVeCSpvcXzfEqbZ7kEgfXf5M9iPE//2G45Y2zecsmTzLd2K9n609jt
elSabHvv2/KthIRQ95Idj/ctG5W4Xy65nKDGn6gm4adyLZrcQDN6sa+LP9j5Ciii
PJ1OEZ2Z4WTLsIyKCVmjy2m30hHybiWEOROZQ4C5/c9d5ye2JvjyC5EMa3/r1ffR
aRz6B5gg6/1Zds95F6BFTJRV2J9w5TxBfsnfsb3Na66IztQDwQCAaI4AgoltFeZK
imxHv1i+ZvY3/PDrYVUvp4DmZVF11KMKxHX/Rbha+LgJ9c6LH4DZfvmUJCKqE0zu
61peoj96v5WZddMEdgtdl0z5yugRXb8CmYZdzJKX5dW6XIhq/+DFfzM0GJlD3YkG
j1d7yD8hDVc0nrbUNmDu72UmztMv4tkj1nAt6twM/stcnonGn6poDJMKtWfp3iTI
1W9XfmiEw4eI25DZjRoZeY/WBHhU0Vzh2zurRGJrHyDs1x61nIwSdVkQS4cx5xFM
Fir+DrJltX7x8WoTp/OQPOmbiaZShqkTLNhCHHE8Pj6fboi4MUMJw67PXUkpCFBO
r5cVygkPXt9GmcYgESKLyKVpecj4u5sewIQGIUhtX3OLVM11Pg/2buvrtpJtWm4H
XvwGqox0pSlI7NlaxdA2vXenWP+aYc44lTCx2PFh+2XF8IoDc3f2ObzL+y+/Cw2q
X1i6Xrbl3J5kGJwM9CgY+COI7WS1iHFxVPeNIEL+v7D0mx8WQMr+9mD5Vltcp1nE
hm+Y4oAuhSqfzo2GF+aZXPpquy4nuDJd0/MB3Wpm6g/abqMiU6FOVThgRSP9ank1
CngdGMsEiFGTSmBekvqNDP3qYi9aVgNt81aSyAKLjGGkMhYCOxHsX7yM12cht5fQ
eEAcnsRNLu3HBxNM27DUsmsSrXW9b7eSvWNgQcnZz7xsdvjBo/SVnJ/1FLVCfSpE
OVbtTmzOjQHqhEwms3eXG2i/EwAiW/ibudP/u/WfYgwTZsV68vLtHfKn1mVIOunS
zv/fVjb7lnp84h/d8s1uj1zRZZ2TywgL32thQ6W6JLMor4/jMlXdl0A1E2zoXjoH
X+Osx3Oxcy/5y5S7tNBuO7kkA3CMQ8KpiCOWrbN1o4GyNKwTi+Vw7bnK8IOTmAEG
GyxWHb/zDWnxmJWKM42e/OUK5bBfkDZ/69PcFANQtPMosx3nfw7+puSlVCYlhHs3
u1MwYg9uIdgpQvTN1k4eWAVUFGAfgM2En5YiNZLUuPgf2qchFCjrwPpYtw1f9req
93rrpb8tu2Wf+5Paelqjcq2F4+jpNYOCFtB3iYP8z+QKdchUCVNg1U8jw33jT6sv
FJKBAZYW4rxTii66KAwAV8rZDnjDOAWEYUJwUtUZz1xd81RZtlOf614fvKpeu+0H
hNGOF8j1mf/eo1iwiUXNIzBAF4M5EynWDgeCexnY2BMzcFQHGuTMuhx17kpdYsgq
seN9ImpYSnzv2XwbZdNx3ZhBUVrSf+XyN03ew4zSHFbkjouNtlKc/8fep/BOEe6Q
qGIyiVYNgdzik7VkUIsSDAN3YxJ5ik1ONeu4DFGNoXibn6mVogBRb2+lDp2dywCi
GxJuUbikm+43bJ0C9qN9Uc7YM6CnkbX2LhxM1oiJm2VElB27W2uzrFlNEvOLj3R6
5sTNkwj+PySsJU3fGZ0iKoXS2gFe7+dMqLQiY0q5j7EOvO0cxivGkJzJ/HdIdKqh
AztJTJP3xFSKUnD+EWdtNMBwklDftXTQhIfmrBUAfvLKafiJHz/Xjs+tnUmDy6eu
DcGpGWUUwetSrnodhiUusqw96o87n9/XsF93GTF5InoYmnx9kIlMHSSQDEzi8o/s
nnS0INUyeIyI+A56oy27qOyTBeETJS9VL3E6FwiUTz4s9Frwaj7tl4bblXkhMj0o
q61Yd2mD8NRF80K2MmMDuLowzoIzJTg0D6XYZDJFaAIWxRBHQn2niOtYEnNvyRaU
W0x2aw1Ch9HGe+QYmMIWYLMME8nJthF9YOUjpIN6BIY+PXwAQWYeHJDZWWwW8t1y
1N7tx5TxfsNM8IDKqmSiFBQLeHSY4cfv2Ev4Ek5MrjqYTGkuZemJiTR/JDoKKNta
vyBCyRDYHK30Cv9reEED9zezaUupQNGs6j8DM8xqGyMVtPvLdBhntzZ58yHXblFi
wf0dHT5E4JlrnfCVT/f9xJf03jMMJR6VWWj4KsF5obNJHWKoeL8pgL6Z3bs2136v
dWI3g3H1AzfFwdm3L/DOJrX8LdBdO76R40Ms9tlu56AtlICpK7PbNueXXfdqKIWK
REt/jOBJaz11MH8tDfqW4rJRjvI2dBm9ADnkOAwPlnsXvzmKSXZJz/rbBfEMu7JL
BXekWfJnP6w800+YteXUbIXoW+Z7cRdAOpuBgPgEtGJFRbUN3QtL8XN4RDAnNq5Q
LoT0RYEQaLfQa/oJ8jRL4Y+z//Rd/HYdXJSWkf64XrJq8ALjRB66JOJo9c28xIGh
3pI7Ink2nDAWX5luWa3BLxmVuApK9F8uz1zm1ZukfPeB2eZVXQUNBdUzf8/TvJvi
IEX1GO61Y8V0/cW0V4s4iceebT6LrCXbFb9EmQgZz1WDD/ywtHThdYuwwS8wMdCn
IsDnsQoBy1SLXXUXASmuGdxTbFEYjIXXnypIczEfDl6fhOG83nIMhhb/2H2Dfwcl
EKJ3S03DhTBWH8CkK9S/iQBE0HDwj4eNqbZKDXsJMqMnJ9pQhG3ahIhVO4DA3fTA
jRONofwiDWSvyNgtJAFdE9qTml1O0JpYO4hSC90cmwnRp/0okroYWWU9IXA5YFtj
syEAs3m7qrkZObkb/NSYScScXKplJQ7pu3nxIDX5CY2yO0EZLfau9DWpgyfCI92/
ddf/wD5biDJqm72ySTh2RQgofgVLeZfiVYUxmZYSPFW60P/ZOEKjYOSDxH9McJXr
AINjCaIo91mvJwmOi+KdfUjH+lH8y/qjBpcfT71B+imrIjrVnwTPKEXtkpaBr1SP
q+ND40RsuvXCz/2nwizYL02FVkuMNYwoL9dq2jEbXZe8jfUbgmuWsu1lRnUycHRc
Bm/PiwS/H8xC/ZekHHeKw7kVOdvoT5PgQ/22tHSv99c7rb57WKRDDzxVqeXwTmjV
3x9u+3Rz6fxVnqqjjQ8i5cvrAmwbWmnODziPU+aykqEFE/vVvZe8SixCf/dGbd2V
0bpVWS43d1P7H5FJl4VbAF/EZ0nGrtBNxkk+Pdws6GPMd7LKDq+9FJAatylF7l+x
768AKLWiA9Nuzgta9jet8emm0LD/hPUZ6oSOIvPiHlP+yDQZdIewm0v5wwtHhW2a
cb+Ftm2dTi1riToMjhd5EcQV4nEcsRGTiJx+lBw3RhPTeiubFgVDzDWLohzoP/D7
N1AoxD0crQe4gz0TQ9Degg8P5Oru5vHjCvBQlhhe8lAImO+7OgXJbCYFK675l++6
LHeLjqOs3R1R8XaV/OXhC24pDxrUJSbDUvM9IIalVG7jDgFO9T79TO800tSApHAR
D0zilVjUytryqZRxHaFmBHXlBvjmM40xFUYdOfyGqdDpyps0RWZhXynkGoG6ubDX
DTjtfuH7dGk1VtdzlqLqjGofZfRUiz07o8DCchP3F7jASkrnyXwM61BEv1ZLL7VU
9XggwDwsjTY/iJmSB6wlscC66VqKewxm7W8I0WpY8KLHsylPOWsRKiRD8EDsVJZJ
HZx4sSqmNvIbMxs+mVfhh93kMNdvDqlbnr+2dxJ9TEwNYrVJ3oOa+nZgGlBdZFNX
5m3Yx5OYyOaaaQo+t68tUoCDEONAy75RG8qLdC2kUVrBZj1fJKLMS8LrFjBroUiJ
iIWKPBDpzIjUbeal+pEU3YsD7TR7UR43XBso81LGCirD+3RDH23W5hGMqKnQDBIG
S7+vV8y5TIQHI6EINv0nD8UE4wdr+qrOJHKRD9mGohP6kKFhjIu3stNbqnddvx6u
T5xAROg5LIqH/tNQb1fXviQiBl5nWSN/kdd83L8rxzv/JGlVfI49yycgh4CU/kg0
8KxRyqrseV1bMoDM8LEkyzxjCpG//Cm/5rr4iPE+BNx1fJl/jt/HOnjmGnaWA+/+
XCGTDD5XdEeRV1vX+PYAh7p0NvVVN7QjmC2/U8CPJ51gK1VCqcTQ0wmR5ZJfOwCs
VXPAKRJ6XcP8z4/OXtd5RNwcoyD3P99N/+rZG8KaaIlZj5gPDJCvFRvYso0gBs0M
WjAb+P/5nSOprIK/Bqq3cmKRDLhQJOjVlXUTQ8fT0p72UFuqraxrKzcEcEa0+hDh
GwSkY9zVYr7K6Vk7Rl/2Cdlz2ZPaxLkGHAOYM0YrYtxJntkizYgZL2OhZs7Iw37R
qOBsP2pDS8EuScGs6ljBj6oJM332JFaJiHqQ/P1y5u2jNtX0sfZFblCUlExyT2+3
+6KrOI4/C0qP9uPNDGMIavC01s4hFfAcsGSy+ceFJPVJEuzT9qL+dfmOdVB62CYV
qnsZgsoakskKfvO6s/2s7+XN1TtK8UosLjsXNFItnnfhv4Xok6mjgGDWB7VfMkqd
NKefhegdE3WxU2H+Zvb0MmhMiZSJfDnztcJbPk6/zTOqTiDYYZREDYFkpGWSwATp
ZQ3OZ5VUmczTFiS1siOxZ6Slnajcj5LV7RUez6NxIGJHV4iMUJSfAAhnBWo86Of3
W3pG8Tx2twgS+VxgvKfacX3Mu3dGmREfHJWbbffvk+jGo3B4OrS8+jWeoLEWjYHT
6zuPPjsMcElh1oYEH30YQZWvFVl8NOkG26lFNUun2VLCVQC/Nq6EoKfb1jmQDBFi
3Jy0Gy3aDwkAA1klQl4oKxlhYqtYpV9JVAJn1mlHd5az43p75WDbrM+8KKCChU01
PuKGaQeNZfnP0emhS+xaEkT4vTAWJWncCb9uIk0w8MjXG4w6dFGxWxtD5sWWGTeO
rJhyFbKGck+wAgTRpe32Cqz9S9SGDwqlvM5KWOLy0r+2VhNZ7+YTSkzxoMuVNHrh
924Ye657enIkqlPgoZckKn50CJD/TMEKOtHwYZtGHFqfe1PBDZOu8Oy57CfpsvbY
t8z47aC25w67QBPcJT73CbsZlx+125dNXx504WMVq9TXzRdNSygvGxAAdrj4Y1n0
Oabrq6g8b6lNvnQB3UHq6f+BxxDJL0dPdlgSAFckxZ1KcOn8lefG2Xsb4Oqp9XuP
su32ZXJv89rKfhWLcua8uWHozKfE+ClU5vQaZrPw0isHrubt2KrnEFXBVxcELq9J
mrsElOm4vKJUnUnU0J0fmp9PD6ctUQRvnoBrQYS5uwZPAKGYlVbdO7QJCg7bYSzj
rKY/TvyHwL9grFoVH+D23w2plV/i28HPSP3zBOT6cB2Q3w0F/iCjOH+nL3sXUQ31
+K/QKOnd8NIayuJSF5mhKfjS9/tT6RgMBUgibyDoIr5WfeKp0DmLIJ2RhdanDiua
mAE4/S2UO+vmFB69fMv65tokBC3d11mq9zeXq728N6z0J6psYrLIabTVka6OJN34
fvaRWK5bOEyvGqnAxtd07DRyRFAfXpBJaD1NvCvg4KtdYBaFYYunr3kF4JA/VCOW
x71kSunWDkenylKvL67haPT1Z7QVYiaeGvrbAoiPEv9MAmx9EOWTVivDHK9fWXpD
0bixXmcSM4qD6ea7G8CLFn2RhC3IBVK86sCD6o89SksBypHE43A7O0TM6ZD4UVT1
yt+8x2g0wKwrdIEb/qfJsQWLyzXn15+gSb81oJk8gACZ3UslthB/OiDgyGxlaRAC
DV/3kiU/wICxUzjS2C4Uca8VRo2Fmg2+EYN6cUmKS1Ad7KJvT1tjSZ0dSvC+pJ4W
ZTWVI4y+EF5ra1I9iI1mjd0sOrBuN+BCboV+Z6iej4XThG4doPpFJX8MRgd3JfmS
qA8EAzumLTuVvOO8oE2PLXgpzPupmcVudeOHG/wiQAAL6GE/JNH2cEMAwEisJmut
IZO40mEcnM7s4rVJIFMin+FBNSsVMLJqKWPNu2c4l2iVgmCV68Hrz7rHyHDQpCCu
Nkzk43TbgQLH54hGKPr7F58gly/I/GugsJpWnKpaqILvCbYJRqVxhZ7tEkyixOJ6
tLsrWoxdf6KnfHuyM0JwVLKfbXhhQ0Lj0Wt/SM7ZPCKLvUJgGpK7nv4nPxA7T+0Q
dETNz9yEmrGVDOSvfPihd5qry1nMMOJWYzNLRI78ZMHniJtlJI13pC06ncY2dY+G
/tdxzbxIYFSNeJeLz5opV0Az/3UELsMFssqKQrJkIIspen8d9mXb4Hxg4d/FsNM3
J9MM9VPFAvEgyApgmPPTaVbgYuzWTMpLz4yPdYrMn+9Az34R8Au3tsb7BLA8w4Ym
3TBmje0qK+czo7jVoYDDIXxO6zK0V0MM/N+81Lp1ur89+G2CVizcLTsvYdJ51PZw
ipMHVC1ycPraLhazSLo1ljlOh2AkGKqqnOjXJY1JzWGOEU8syrEQXz5Vnu1YPNtS
EGd3jQe66aFRcfT6S26g86cc1sHqiwzoVl+CJihkzRojDuo+Gi3sxld0CYO55fc5
2Q7u44rl74R5bA1XlzA7kpK9I89qzMWALYlw8Lty/xmSCVqjy+hO/jOLFmEp7OKw
N/ELdIu2mpAyTCVaAS0JQ7owhFZzurRmAquVWMwSRemZPXG0tGIjB0mftj338qsJ
QTP7BZMAB3LEVtGOGj8naDyT26TNnfDinEuVtNgh2UgFUNX0B1HZRT8BEca2u/om
jpP4V9wvc/9moZzMUdTEQ0UrOHpXl7shWA4b6BmM8gwvlf0ADXauhW5y7AJJu5Fk
56U0qbp0HQYbi0mBS2L50DFwq0gepAbnqYyf+EKHR7Brw7Z1bu2keK8jl/42h2ky
U+gVWrSQzpzUjzHCPJ4bPHeKhyw3ruLmvNCRZZjj8wwmgA+ZaX9MTS8dj7Qpqav2
WU+zY2+Y+tlX9QBQ9sWIuTqGeDwusZtgvYAn6c8+hHlQOD11f0CieUUpOd1BAnjd
VGSBiOYq4ovSyNhruItLHXSmSroXMIJ7x/zLOUEOp5l3gI7azNcWd+1IzPztxpmf
MK7kAdvzYwghw+4of9ohZwCegqmzcGq7TFaIJImO+fPcsCVHy42uleE6hhMUD7tZ
yxUK1zrZNbjTs7sTyNyzar4ekQlmlurX3lfEPOs4Y6JZrW/BMXWE+LkHG7DmuMW3
m9qskuj7vyLncpsW5mi35JrOmv0IwCDtdZ7aATzpNDIqIOkdIKkF7HgK/6cCd7jP
ckdZnfBOBucGyyNb5AtrUvl2M+Ddu1oH9wlICqmC0XurFnyGmaOvvvVpqXWvaH0m
cAJBG+rmfvAsJIyQrAYRsmcgcCT89oKJ4v88jcHqZChZe9Jy2lo6i70fbo30fOQe
XGykYHF5MSaS8f7Wm/nJ1G46ilGmcltXtz6RU2AJM597rYEOr1+Rgrw3yaIyP4xe
Z0Ewm608WeRzn49OWO+s254+RLa+LR6aC6zxcf9uBIdARhmoO1xgIFi0jhqSY0Pj
mQkyHfIzL1GRt+cAy25xXTS07wCOOvv2ObEtlMu9A57TEo5WXlMXNz27wueVnlqJ
YP8GMe5n04rTP3wyvNZjIYRiK9DdpR5xXZ5x0WyriP254rMbUdT1LtSEYt/ov5Wi
e7ey7vUwxHn+PFbj8+sWBvL93Y9JFAJmnltmhL4bl+GA5RpEPE1glMux8MRzfMBy
OVkoAShmNC33KGa8nQucx7IzJn/q1wnqxHVkTJNesxSzwm9/Xc+Ntjtv1eSqN27W
PB071C4zxeph5UGdu3PjG1qygu/bAc6vnr2UHKeZTuwLGlBamUNPQn1KwyVGm+3r
ob0+mIP6oU6WhZ7pOPeGoUex4EMF71GgYIrFkzTeyrsZoYVjW1968xehSQwgyPlf
AIysiO0qXw9cZTedJ93upMy+Dl7sIOXB/9mDT1xEa0ZYVv8Rdi03SChUgG9/J6Eb
smayV1rOBT9o6r9fRxDrW6RVWNcEKNrR3JKp7uMUyLgqundYrRjp9aL478qzOdga
NohYnfBHPTUapkvvbktAgci4XSbxA00H29yTswCxfHnlZH4z3IR06tRYhgM9JiIP
v8uNUOMVVFdluIH/JXu9eMnKk/fMmq+YKSCQ83VRVydHSD5Oqll1L9dXXUgeRrX2
UKr//8mtXwzB+hnKiek9DrTdcZA7FRpzjQO4HEY3EZFj+TLkhB5mEBYgOYSW7V+k
wmqjqldDOLM1Kou4zZd64vEVv1WGcU9T/3DLqNjkIbT31hC3PRCxl2w0pXQNQEWI
WatUcXw54IHUCTDwyxTyhPu7Tx5g4x7+Tk8tTLjb9ngh7fpypTpX75iZLFnafQTX
MTeqAsMvjJQnbnN9wC3a9IYbgAVmZC5+anb/SUW8Iyt54mAUDIeebJNwZPumnGN6
qO/YIpZpXpLH5nzQ4uezTaU+d+j8X0L5O9DQLkrSbv7LRmh5yanvtXPg7i0bmsVN
JgyNXYWtZjFUG7rXlEy4uS2kqBaBZr0B3K5mGEGDCWZ2S0//OF/KNOvfir/HzopQ
+9WH3hHSEYjDnjokE4U0YjhIBvOc7zLUUhCJdNU5sVeqhv1nHBXLYA+765EU2v4Y
JvRhYsnIV1wP6BMK63GpWmhfR6J2HqUNdrrx+0si9SZYkM61dK9QfMF5LDh88nAk
y+2IFTA4yyIcvh9Xx57InHgnjZAct02ebSsJ5FFIx4/pwVLSVEUCn8XJdYIIcu4Z
yTSXieF1a6ADkE3/Re883lIYVis+QNbAZfx3HAEhQX6goUFNM4FvBEv0kSz6+fZ4
reMnpYva67Q1C/JRpn0eeWy6QGlQB/4xWHAEw2kPmp85LdZ4tkyE/6V3Cun58tZO
ovfwUmhYq8dGNqEQ8/WjbD6QZaP79OB9agEPYJal8b5wHw8Utu0PJ8xGTOW5C6im
YxrNR47o+RUHu1On+x1iqvQpsIWOpDUbAsA9/iAPog3gq6gYk7EojU8RWeNliGdR
ciTD8U7uxApflWuXTJIgmqK9gMQRj6Yz53gBCjgPLHJ7WqzwE/FvL8F5mICz6Lr1
F299uaLoGpgPw5WaYj1EbFZGPWyoIgkDEi1XpGRKW72b84vHbsoF1ZmKedPYnNr+
Lo3IGu6RTFp0nrPtzBE+dpOV7E1M8D4PqtZZDMzf+G46qtQ2nZDlUBIp6igZ0iHt
BMX+Z8zfzN5GA9ZRPbuzc4x++hU3AnzxpvDfiJjkO4/DTgfMbj7X2eeDlp4EK3A0
Nke6z8csBgjPpRkkbTSeiI3c4nQ5wydLX+BPQrOA6n/x5BtJ810elBih1hi/nrQB
82kHEecsoZsX35Uey0rQGIOeQt/Ki7QqOrEhRbOAcf95XJW5qA7BlhOu9zRBPSXb
+9s4qyQBJpOApG7z3o1ialQxEGg1JdWTN6DeT9U/EkeWz6RBwBzqGJ1icpfVPEMG
kv9bnrfsUWBYSe/Kyn3o0S74fEMzuGR26KgJdtieENIRAwpcdfuR3yMQmJpyrWhh
JkzSCAw/duCOUiBQoSWmqk21rPFi6MxeGqYLvB5aA1Sl3wQv81Br5/VRoLr3fIO0
qNBxNYHRWuh25q5WSGZZ179WzCS480s9joiVpEtes1EMqsludTjWj7pJBDE4ekm8
MVkK6XuRiCdYY1CdRKqSlJjq72S+gIqET28UysiVKRDhzD5qsZLOPTWX8weVLRgb
sfbBwPqFzRjkC58DQilIOdYigLt3veAu6fiZ84xYTrylElnoeGqfWUNrqjAKwcfA
B+6ZiPjXtYFkrAcZIsRzF76Kcc2eCkO2Gm9HL7BZjK8w4pQ7+UUc2TNagDbQKin8
ISMbHxGaMygKznK66riOKcnBSPoZhaWOXihMV/cdR9FW6O0NLqu0BWisMVAexHYH
gHBxaTgkLX5o/jf4LijbYE7FdBGq8781WcNg729LHEXBbRM+bP0tdqbAefKGOpPF
3CdnNqztjuj8qSsygMnLOBN4gZFfErxyE1KWroQVmK/66NA8Qk5okAI8d4mOO9sK
7UxCmdoAnIelavzTlQeZ3+eDu8ts9seT2z7twIJVaxy+v2fCeoW+7eHDvPUqbnKt
cpF7GmrFyTLN7Xsr9an3fCxH8WQh7SVllLZsJx3lWyDqLogicz4jxbj0Yt9LFq2O
/ubcC8/X9K4K1b/vKMuj4mpKlBwqfGKtJ/oz5UK7iSls4mZIjQD6AUy9WpX54DQA
+HTw8Dx6gvwPLH+dHTpkVYaGIiOoxuyMama5ZVwFyfCj7OPUruH37vubBkQhFcWX
/P9p7omIkM5+9y5cIkFbJRdU841lGzOBSQ6T7r0dSrj4BqP8SmjBMJKLKLWqMLBD
TjBnGEhK7tYyF5UDGgkx75RPwEjtT4ITorWAn4UDC/roztxT8wk1AwgZX3N1Ar0J
u8Dbi9HEH+xSdxUnBNkE+0IfdDUrSPIvE8oiqjH/fhE150xcHCRc2Vg4FtXYnoUm
VJcCryYo70xkrYBZCVyxotI9SLi5RfAiwXScDnY8lE9CBjHTjJf0hLOvuxIQZbf3
y/yjKKQOX/KwzRo6q/SxpWJ7dPe0o0e+uOnaej4PvkOOkaYohH7ut5IooJ8EPba4
fzCDZ9pUE4DBvDijtZZngLfpowsPzJd8WzSQMrSeYvBigayyxe3xNSS6d7HeqpPD
zHEUsm7o0CQWdq/MO8wIsFIIP3Pd/OdUpU+fWrqXYwnx93C6j7aod5xhhUWtCDw4
rZ0yUo3ymds/MaXbA0XleD1KEm/bBWKhem5p0Mg3BB7Gwz/T+wSDxDH95wlrdwP7
Yt6dlOB26DEmM8RuXFS8snGxeJkou9g+K2XkYSkAksN3Xx5US7s2suTlDY6DADII
bgbfujCMwHMflAtZeV3zRHyGToERz8PRPQWp8gYDZwh2EjIMN2AAJfpxY4xpZapD
oOVVGnUTXDSQreTxUjpFc8nlNui4EWYQpfmyOs21LKREUZz9OY1R9ixOJK1n+01L
pi+zvaMjuqbdnGmyKBJQzSmBUjGpp0/KpsxuCaa9YhxS267zX5zuMBcyJpG6cjjv
DgSNKl+OvRxShmjIpHQDXKgcsddrBqmIlGFz8Its4vhy9Dglg8JRv95Uuumiyk5Z
Ft2FLIWgHEpDGKucGQSl3wB2ACI7c76n6l1vZiCK5ucHFdH5wHJY2oT8p9TwaWdH
DxAxA/sLBGKUvQfYxJrkJ1WJ/wcrjhJ4f6hw9AKbnQGcdBGZvI6CZpvF+XKJIA1J
AtK5BeVaxdDNqjV225A6n4IvdLx7rJNcuGkV+ri1RSo0wHWObQqlkiOKllW4GeW8
7G007XQQPvkKru6GHu7MuWNuiJ1WW9M2a+FeaHJPB5TTDssYAJRLeCVUuYknBjoQ
8gp8fEbq9ugW0nOZQ63UvE26M2ceWRDW7e3MnISbvmRrc6Dnmu6ap0ZzWE4a7ITX
rO2l47XYPVrQNGTSaG7Of1HXP6X0Seg8bIp3KJiSmMYlNNXKyKP+K2xkd4D+AZqb
Y7/42KJCIo6zwgPHqJrdQtSAor+mas5vEV+qjChoLhjhwc28TT3/KqQmD4Y9jRcs
YsbQcd3pn6JLT4duxdt0WozJWS0VbkqwdjTqZ/irOj76b1wArEEDzIou3zCosUFW
P/oIvSa2C0s+RVgN8Oq8xOUj81LnFafDTbkk1dOFdSYXENV87Q5a7ubMmf1op7cz
a97yxNl57316hUwFHoLDW07dFHoxxoZRRHsyG4kWFUyqgGTlOvMtyvamdmqqWnDw
vgyGeiVEhkbyokiXa4AOhcUfEIGvlrplfKKIWBoRNo0Q+qYIkrJmY8GyIO2Nm+ft
Qm+cFV6IzgfoyjpL4Dt54slRgWdn88Awxc6FxxARp21eQIgj4zfz/darl/WYZ4Fs
BvG/BQNSifj+zHCANU/pxgEsGaGeRBZDlrPp1cpTiIeHeLCJcmJzyexNaWApYlzl
2IdkjYeKQEACoacM0AJzthjcbk7ONGyuyZ2GBQN3bzhvGWD+HYIX+ehckhYud+hb
/bhocSuVLh/oWEMLRcyOsaEAE1g4+lXw++2sUySXh0GAUPSUsoTCOYpH1KXdTC3z
HCJzNHh6Ox7EK8B2lCAR3e6F/szUc2SSmCV7NLntpo1pyJ9gGkTsypKC/aUoGqCu
lHTrPCLrhRnp3CQyCY+VUbaKeWhNMtZ1pwIHkDecLLhJcnVLud+XbO9hgHpcfim5
4aMtgajXUMiDezJyxgSrmQjiYHz16AUXuRFD0WgtX6u681VBHpT1z5C3qR/ESed8
LImp95sOxGuG+Rgqcp6F/1S/1B5Z5ru+C4w/NJ+R96k9N1Hk3S2r0zYdL1OKnZnF
00YlIDJw8eW7+mIDfjr9dofcneAJiniSclAz4MYGSXdUmmBRo0L2nlGDr12bmAOC
zV73rFLmulYxLLrkwnHHPdSZR1q7HfoBO1YCYBoB1tT+SbHgYOIgbcXsLCNVzn8u
EEL4QrlgR3/fvIiBVuY/vsto66BV5ZAZxL5RzyLZnK7RLxTKF49FliPVyIB2T3Qz
aSHE9YRSc/etXezdyeZ6FS3UbOgC+YxBlJbEkdPVxLPzAXKYy02xsSCg9qY503Om
QDnrMbZmfCsYkDYzCkF/0XpRlgHPfFAKh1m7wUHWYjjF4XlItwXlP1MzZ2vBWApr
Bx7oxatbINtl5KVSmdDhOWRqzjHO0lL4aiFKlpJOQgxvVxFP6KDXBFM1k5lUSHlx
J0Olubdd6dT4VfV3Kh+vHWwCMF9nqgY/9VprhH8eXJzSTf1NexApVftdU7RPkoKu
tXdHwQgNPb0Qti78rzke9zoHhG+ATrsYcD7+ELti+xm9/jR+g3G2/R8ggqzdBzrz
kbI8RSU8qsOINPAwPZ3GmojsxA/SzPaCQE7kmje3l2KhiYo1gy7u6Kn9ci32hW3p
ZyOu/DttmT7BhL4v3D1CJkpO517DpeFSdYJ15nR3lU9c5os6QV+dOypF/uS0RkZZ
OzXQ0Mx4G/3HjEoUnAi2N5WvBsiixFxGzdeOwGrxwA6FMhYTBcURL5H65ykQAL1q
ttUEC6ZgUeA/6OTJoiM2O7HG+oQA3WOH7ZtvrQezIYcvF44q/fKhNkJHQ/SbrrWo
rVKIDA6fztTBICIBtSckurydOoFSoLtMynRwXWM9IWmJnL10jduT5WUuaEcnw/vu
wiqIASWEhjxBEj09nMkPnVlREE9xY17s0kzCBN1W1/ZQ83USQseJqK0AOwNjJnOR
DT9ikxWSn09l6YsRDW/Mtt0scxYUEmtaMa02TBJiFKKDe2YZKORqY7r2IKI1JTuc
2FOYIAZrtrNhEKs3Jv2xVcipR3eU6hDLc4CoLZ/+n8fHVKDnFqUwk7U9v61x1hOf
oQ01Xykm8ZhJb32kLMx1tFnPaRDQ4CBLXkRezQFoZzqG3ZiIWloQG7SS/L05ldK4
d+mUBc+agn+Z+q3CiwFPQ5ZZweHPVCBzSrrHK4MLuRnQUduU5aj8rkD/6umT18It
0PYNchzAOGqeV9S6xwPrVWD72TyTNYR7B9NJyomz11vBnwOPKeAz0sukMT8TEzyE
j2fNEevf6p3IEF0oYJXOIirPnLBIa+JkNn7sb+FrtnEoLTLckAqVt5Ua0Fxlrhz7
snZVxs173JMt1O3jGdKg2+MHyusihkqQprMAUgEpyoCND0WOX1DGuOisRubrUABg
vW1VQoWK5HfimnbJ8oGw81e1ghUpipSKGAa0JUfsCk6vrOVly7rgxhp1CXzuVGn7
ye7rPO0gJsPl99wy5VG0oI2jmbwOahHCvfDI9Puz/j+ic/DIepfZXXQZTQGWRibA
MwPsWr/jFWOLmuK3fdGG/98yd86bzJW4Vm2NcxmhA45CWiz1EYI0h7auC3LiKY/K
ckBSKNF8v7kXEnNCokBDbNzkted9LpJkhr5YOcU3uZ48+ZREjnrndUMmopo7YcPO
meI4K/XafSAeRxfg7mnUzozwUJOLVoHFSxU027d+7YFhwYdAxRmgOLTI6vIMlnCb
78rGIssZ5VgEwF4QRRcocVqicPF4iHNBDEjTD1yFCls8I37HiR+GM/IY5SnMja9h
0YXzYociiqbmu5USw4nWjJHrFQj6lNbFVvfo7JdyfsYhRyA1FEknHJQC88Xxq6O2
yHswAaQfSeQ5aClMH3Q43+gBTR+Al2DQiVvCzX0B5OullDa/SkIa+5e/0xufkqrD
N/IDr6eoKE1Z5zEwnqIb+5mCLfyYP+uKuNfBoF3c+9bk1eNHyu05rSyL2UMZjgtA
d/hu1sCZwnqsYDLJ1e60d5yjvvqFvIn92Yp36lLYYjWDpH2cV6xJXf6HdDTpU/BK
90ypA858Zz1UyentlaP1ZVdcMQ51CYIdcNDlVwzSGdIlTnIZ1v2Anu2Qhz7TyPFJ
zTg9ypeCAcM/VCd3PxChNaClLltcuvnekVj6XLsl4/hbHUDNUusLfSUHNmiMdEy0
ugtntuDi8MbNOpzynX7A+Vsm60eZAf6AO34NOcJrtr6jDQoqYcHPc2QDcZyIIjJt
sUZGrqIvrHE0Nbhha4OxNczEqvHQzPlTk0QvzPAD6yxrimL3se6qzXUVJ8/ySA0B
NKQz7gWYd9Lvwy9bj/7ogeFEZeS6rUsD7dnQvOz/pnnjNcbDnS2/f2y21byAP2rH
4BtDnwT+Ml/DNKThgrCMLfAWrVBliHb8tbvIcmv2FYrwlEfMnCBSpwsMP7NL1jVq
eNSzpnDABtba4ucotrDBDURRtf224qwwjQOcIqsS1mItZsBjfmC7oqAbig61P/jz
d0EssHvgXsXiIF2zT4L2adOBAF/kUlCtL3yTJO/DESa4oJCoFcbV2XMRYUzAiQ7n
JZbU7dAWyisBwh5UvlY07JQDPUgnwT6M/0BfrlrkFaVTnatRpcR3RRU4pQ76BLyu
6hIpSoDePwUP8yyPypAtRwTcUuvRZd0HYhBKpCj0iPRl0yERLLIU5j9475Np4YRi
5AIZaoJ5ZV3GOy9gysfjxCHCFZ18XVn7zrKJPKz357l1RFO+aL8oCaP4omZNA/vM
AqjnoG3w5JcvUL64wRNBs3xbehH0t64zTPZ+AdMBfOZky2bygbBv6sL9rpg0qpiv
HfVCTqeyqOXtS+LzN9JU0ii/juv6PRDtofKgUfYBNDYJ9SOzwFd+A5gjEfNXVOUS
1q6IFDNAz71nEm/oMxE6HT9zIKXnWrO1TED0+Zg+O4oL1/Le1vJ5/FtokwVBn5k8
K/DFTOBDaVbL/0C5bvUW3NgIOeKQwblUebjwV7mv84gnLinPQ2vuxDOvRRCckh65
TcT6rob35Jn/rLiNlsiZKhRtjVzyzMGk03oY6e9oHgMoKwlXA8N7rQxAfEV/UJwy
rem4ORw2pTH2Ux8pdinD5NUdCCNos3YyMcqegWquJodPc9Hp3CaVFpgtzvZW9OlC
/P599cuTfYJI8Bge6lqKVDybiJy3wlmFmW/xFb2V+vaH0mgpe1Dv6rIfGVzHC9cR
NNFBw7F6GyLYPkUaV1heNdCORjDdZtFYVDhg7bGw/g6vPRQ2B3S01DTB19f66M38
Bq74mcfSDiDnRgSek6h8t7mzPAc6KIfrBLFqh5gV6/JayN6AQ/hfv+uf3sx9xg4O
kpKgV05mCNovi2VHhQ8hdasoxFX9uENBe0aSbVVFgxXVYcFUfML98s4VtDKSEa9m
ozTGH31R+q5J9DG2bpjdEeZCgh6NgQNR4Oaiit/zz/xeKLEsDFLPH22CHiPVUAPF
Gd8G5igyBi11FKTChRL7RZJpI2CNAmyk/92g+8FPTbrb0AJdktl7XbVEebERZqNi
oGblpfF3hxBpl+HBmnMkcx+RGdyLL91wqYcQGNXEnAybQTLRhJQYd/Nin6Ewyo+n
IPvorV2xEGK2fXShPivxll5J0G17dWl666RTnJjG4PrZ2sHKa/qcp2bjxaJ5E9gu
mb+rnIraF05JfuP1WMaE/lPK2JpDwpPzjUUZMWFAMKqAa744f+RjliGm0qyMRgDk
OMMrwkMFgEiqzKOSF3SJfzk6jY1TEQGZLxqRI4fSpRVKoT9D90g3bfmYsA2sPeKa
cgOs/Pa0Ctu94XafmQtyIHruCbBkYmnvGxF1RjZKDohMAHlpsev641G/VECpZATc
fr9Ftl6bsNTTKmsOWYgXOESeT/hF/FWt+6GqemIBAVz3n7uT9bOG9ZHzdu1V7bgN
bgCCLly7JDSPiHeKC6gGqTVOVM8mNzZ6pJ0+pg9gUk+PjfW7BCSH8De9L9QG+c3H
sQcnb0iMOlGRiTtWANTNmkyjF4GCqaKZLxfvGnHAsZDO6ylQdyeiQGA2O+bPFqnU
AZXqfbL/D9d+7dKNPUMeO5PcKSKcZ5Crlheu7+I0j5v4BqA8PM3HHoG9MWa8BXeF
Yulq8lhf0sx9nMqm9oL0InQU8KiQ1N0volLR6lMEdFv3CEnfT+Ou8MsPKTJ66kHa
NXRHzOQM2HPDJoNWxL/7FA7XzHYHIX2jCxFYpdMz+yTnT9FWOkYKxdDQrmd2xtxF
E+greyPx+71U03Rim0bhB33ZoWRGvUQ9Gghk3NsBrb1vSgWQlPutSbCcdxDdzOES
tJThNhna0whFx+yh7EleAdhzbIMJpU82bw3bQT7OqkbuhZPO3dZvmxqbwQAFV5oL
mCxaHglZGESJr9cEM+iujPQcr6wQfDLcEF48BGAJLy4FIUFG7XZ7Nc9M6VhfA/xQ
1O4+lJ7Vp/pqMJebm3xK4hjOo6AgceTAa4YIG/SDdCprBIVWevL9XBEY+ckagwCg
FIF7vjCb9Ho73bVsh0VzMJ8RzzotQpCVwFNLe3d4y2P7IF4zTkE5fAjqOQXANCRq
3EJ8ZLiSE8iX5ZwJ1+eW0qRLzE2Crpxxzy14CF9Tdy45tauMp4V1y00Gx+0jVsA0
aFfBa1CDRJiAAZl1SH8czcOBSoD9uuOYc09mWmXTa+9tBVFgGgXp1TWBBpnhVDt3
dSu/3Dh6A3oIf3Rqd5GUI+al9MBljQHXchjwqpJo4Ljipo+rdT+aLfPVYrBfALLo
3oXG/RbmGEB8DMsryaC8t7Q8o31i1mnfpq3ZMy2zeBQJa5mGsXmWMnz7e91SLF4R
DqSx46rJyzNiBn+3FrmAyQlRmCjOrcUp629N5Z3tHQTXcm8/7lQe9GYPzCQyT4DI
6zvVhA0Ed3drIgVfiA1ASm1KigudR/fdel8BskAu4g5uzoAg1OxQ8KyURSyatRwp
g5i0/CqItA+Z1O0VbP0HRwvNLWg/haEVxJlj34rBf2M0nSnfwIsmdXl9FQA2kIBl
4efafm/R16izah6CyIB9qawqeG0R8D8rMQBFkaRk2yGs4jHhe/6bVjH2DxPYweOR
tNpJNFBLXlEOCD1mVDagWvwCs/sdFzgb21gMjvsyxN1LFUpNuJMH/zcCjEeq36tl
bQglOt6pRJ4foou7P45wv7Ooma8irnmSX9VAuXYB4F71hNGyQWgTqwSPGngb1+eh
O07gd/0RpceYEdmGzzCuFxkPvlwkg650zwPNFACd0ma5hMMYzjEL4pLxVrpiH2+8
SF+5tffh+xfjt9IHwzhDfB4uvecfGcQFt9U2za0m5x6k0SPfa+MIJmqVGdEUii6v
xBsBfXGxwl+JHvFUkj8ICAxzoOLJzcNCINlJVqhurbotvD5t+9bmgoSJL/2gM/47
P+uoyZ4akWjqI7lAN1wfS2XC/h+IcF9BY2D/Rgz5JPXX6yWvl5+Fcmjgs8xq85Lm
ezJxJTV3DRxar7ioNRpmf7eUz8Evohws+k3nX4DuYRvFOFNDc8WNhwDn7hRCyrv9
oV7wQQRXqJfom2mG+tQUODEsPrVQQVxNSQGDHf3+3a7Tw/vdyUzb14mokC/BWszg
bSzXwVMKDHqoYtNBE+QY1ofubcz+yVwD0QTuqm1UtMuaZ4q4dS1lSDyTQlaUhbFp
SngUQRJUjDUVlYBlv32mvfvKARRsWLWPT5smIFBIzRKZuKkS2Ef68l/ABMS6Y38T
EUPawArCGR9n2Q4S+a2+xdP/OdK4QWzfWuzUkgmbYdsvbrHTo7UfeMPtr8tAzllE
9xFIXpmlgL09qxPqg/HONa6KTcQW/5j7blFt/oQ9i4aPAKVn2QId8g3x6keV78B6
kzlv1f1z8O+weVW0Ux0zSackudW7DOydVcbhWVzDr1m0msrO32nGQwPyH08L0Qcq
fednEHmkXnJ6+dVDoZEjXw0mX7ugknTGNeg4hWPwoSLSOEUFCkeNaUQgCI6mHTE3
KUl/2ozd3oAIM9qCW4/0Tgru/HIFwg7LUoTO196QkzPMYGRJdAMWBC6k6ujsotLC
ivon5E9b05H+DNgps0zjqqyGkQ7BQC4iQA0f0kBNlSQHqz7jQbheiIf6J+2hx/Q9
sGTVJPAaYis4h5tfrGxz4pxP8ErgQNxN0mh2Sr5dJPCF49aCa5VBRMYmx+ObyDyc
J9FxL+hhlzdDy8hgy/WzON/XiQ+63daSorhhtLCP3b9q6FNIVUpQBBFJhif9U+gT
Mfv5ToHzILvMsNThOQUbV7K/4cahdqSVy7myyC/RuYIW4Ou6rBmTiua0PVPc7Y1z
kQq/UPnj97VlzsMEidMukSwZXE+GsB/NhrV4vtCxdJqL/bGZVq7lvfesooTS7qcU
d5FbImg8G3qvV7g8ap2dDohKUAR1R7vbLKXEBjY1adj6/NymS7OCWkLQ9Vno/S1o
Wvogd6OdoJMozjAP5L8jSsCQpmiqgOND6PNaeZQd1iJrA3ctBby567OK615opyp9
gdV8ZwtYMOUf8MF4Z+WeRNoMkSXXqF1x5AbPUx5Jr2eumhB5kr3//ZG7geD3unck
etxa3gzePe3b/rLjwW1H/F1M32aoveuC+mMOKhFHI4bDQXusNoX1amiaaCSU31px
Prqm2wORvPi9B9s6Rc6HMjKM4DTOfVL2QWNwXOOj9GcZYHiKRr5iYRkzk5eo+xd7
VBwF90YENyidtqyi18dn/49shOdWIU71vr5DvvLYQjv3IcIIIKeyerw3Ek6kZ4tF
HvZig+4VnKYgeILU5svo+F9YAteNZADbwpNbbZb5HH/fiw3c4KcVItBcNf8IEQAg
R3UoTHvxExMx7/+MV/0LhHNgGKkbK+yF+hU99Xr8kNu0D2heNksnuek9mRQh9DuW
zam/GESjOflYNVDfphqcNdGz1Pl9fVZ5zq8WFyUOmO5c8n5oCRSQc9NwNeI/TIaR
K0qyBl0gVdVrYdoQiKrIM60yVXv44fp3ThbGxoSmcI46zlX2N1crVeY/vKqrzbgR
56Sqc7bUxjtDRIr3M8HsSeZi5Mywh4Y8YImWlTVJ6KOeRsE4ENULSqXnmBFVwb18
XCr8pktnNWSEXNE/4YdUw0YchjDJocTYVaMxDr0+2/S6XzkDJv086BnQjDBWb0TE
4rZFGhh0AiEFfrXbxh431IAkywZrw7lZh8aoSjcnIP5uPTOo6uCiCEU2S/PUEH6j
aaBp4yU9OQiRsX+xa1MDGmoK/oevGyRfdiqL+Ts9MuWNEKkRo6HO2gnaSqT8e6AR
/ikrlE0a/M19vZfTz4naO5QHC/kITtqUnIbP+JWxO32TGukheAkxhHZ7Nv+T1jJ+
FUtDBujWT6ZgYTgQ23RE4ftCEGZpc5MOqcC3y7jAZhgFsgC1IWUcO5Njx2knTymj
wWMTdzVRUnqtkj1mfynV8/mBckrH8UdV52mE6DgfPMTh9W84U8v9i9S9q6cl6OwN
S92olH1l4ltqivoi2bZQz7yufBXUIaFzZezBHC06zTsloiBMokLCGS2OXTemXlol
R7PHHnyqUgXaEU8ricu7p1TVT3zhuO3lYEMyO29MDIGcmyUGJQZTBOqmrh7syaJs
itfmM+dS65cvPekDfq8gNtOyR80B0fLpQOEvsq3rOZbiMDouVXHSMYM+lY1YuIlE
ijx07gIff0XBVeJagvYICrwPuw6wZ/5RmHz9cavlrzSisY7Sr7hSQ4k/yPGeZj9T
fODozb7lThY0Cc796XR1ZWov594fTzfZ6Jle5gFRRTyWpWj3qH4RXN7QQKlUktUL
gZBc6Gj2fakQyx4SL9XEbF5asgqbJZZoG4G0RLfgTtggXODJt7iQpMOMLIZm/uC2
itock5ajSesWlczde3S3sU1jm//rKXRNZdm3d3pA9/dSdrt8czTgyphcb3Qovwsg
vAHjjQPVDWcrZpHrjJkhS4PTaErNrd8lCmDOhK41Aei5GSB9tKpVwwOpvtxjJ0GI
UxdH40tfnbexwsPh/7CAiiyltWAAjXtKbjhRcyncTwq3uE/uGZPbICiwLdeE1xhB
efZkALyPqTTb+z29pCRKzunYJ8IG63FC2mbX+V9YdLmyJWq8SwsUuy8Fegzd/KyJ
YMjx29HJQbOuXq+h0RIV8APjtBAtlckDZwrvNp2m9P7BGrLln4Zm4bfwprRDwXVz
LjFsuajth+NugUfrQGts2+txtqjDM44J/QdKlzYrbGp9zcmrpwa2EkKCL9la5cC0
RV2zq1Q/gcuk1/G8zgflXtc4aSdMqqQXhtIuNhaT++khdcEtCnQdF0qL6Ot4PHD3
d9EWs/ROi3dBFzz0Naulgn54ESMUL856lB3AFT/3R8aIo0BkXshr2DSmdRfKYHWH
05iaFCGfMpYF/LBvfKFl261JYNGu5463/oOKbzWlJ5M+NcO515EqWzBc/LzMMVzZ
GFUHvhWQeWW03VNvoJKk72fwHx7ftrsO+Y3ejq23coM/xhCDuB26hyxKA51fNm8Z
tQU+DzsQq3tLeLx2TrwWZlftgI1VkHtfwbVSckWLzxJSbLpykv8B7sBD8ag0pueK
MH3TYvl71RwX+pqFLtPJX0SNhuvqiEEEN8xyIUXfIZzWI3YZolTytoDPGOEcwdMH
jHBJH6+eKrky8eOQk5nH+hPeRk5keBiTkNbvll0nf76aaa3qW/Z1I7G7H765aVqZ
TQqsofKWYom7PzVkRhBLpSbFt8ATn/+qUM8Wif3stT08ZiC/XDFyhGz+QdHbeJ0K
v85DzRL1/oXUxeUsEk4fPpJ617GP1GhTNZ0kInfij27vwNPH+o5h2MR59B3wAXCS
Hc8ZUYlLIOUENEkww+vhywzvBQkxH+K1mZFVrnCMF1Ssl0y2z+DN/zihOMVyL8Hy
bY36jpnJnvbWEGXU7OHlhpodAERtCSluwmUmI0Yz5ayT4KrXoSjWA4TYPDYQT1f0
ZPSmhJRlAK4ZJWfXXjYhJIxkhkDPS+6ybiy7p7esJxP1Uasewm7IU/Xt95uHy1Go
xSNfS55hDdnDYz0hBo8CgX4ADn7ZqYD9MWevRnQ83EzqgKIc0lyj3MIpT6wp619a
Bff6iedVtLKojoC2IUC9gNSSyDfMlC6uaZ09nzjLiPj1QpuJVoFPCBdULYnbIMOV
T5rnBzKXWWsDlPbXCedD2uLkei3BoMfH9yYuNAoBnZjO7BqvsjBwxBNvkEf5WM8l
7Tf42fJQYYy2tUB37TRI07UrkJ4mMX7/OkD+Dr74zZW5k0toHxNsfg+nvOPjAJ6/
qVGCUSvUn9/gebwoPUb+xrkqnLvaHF7kvTHrjZ67Ke5jKGgqBuPcVGWRi/tX3Amy
D8EDizcuWmoJMDzdR/LSeYv+d0w90YULLxgWWAYJdu8yWC1ko/kydsejx9ZhW2Xw
XGRhx5U2X+NvJJ4VuOdJJ+kuMqEg2BHf0hODfb8TIav3pEAwzwlrIxhzgDZrb+n+
c4RTSXGc9fMgO6SFKoVUCCQQKvZp/bZAuOqyaqVUFV+NXQsJ+LS8cN2WlVqaVv8F
VdgoZnnyNF6znJ/9BoXqFpdNE6QzETegClvbTVpwENgBmEPQyDhjYR9UTzww9whd
YRDyV1qqJjKVMjWrxOhOzwfURQ1/T3UAwHlWzEYlcLmoQsh2GI88KVHrXhLZVMSI
XQRJBYTxFe0w9e4yEqVnZcPWBIAnebFZ4zLFQf7c6kHuxKbiF34b/6isio2EbQvb
KHvFVBT8cxYKrx3lEhct/CyGAqM3pdlT+zVHOhMLvXmhHlJHwGstFkkfAltO9u7q
5kSaruEXpRVWIjOSag9tBQghq30RtQQCLuYSBhW8s37pJtlzP4Fk/Dy2hmIObJf7
w0LhkO5Qvp5W4rDkLUhvDsGijoYdGi8BuGYksFMZUCiavPoZ880Scp1pdaoRz0ML
MKoacFjgsk1V7HklVCLjgMWj+FFNU/eB3jC0fFOhwOZoO88ZfNoJc9+BK67TSa7B
yJYCS9odMppRtPlm+eQ6jNXULiwUjMD2m2Pz5yIx+UZ0dNEBh0XP6IF3B9GgmH8p
SiwEXWUaD3tagr/ggT5RVAkXUoLNHhQHY6/w2NrfKDxwrguYKCsVtzXwLUbndsw6
titvH1NM7qbaT7vlVWqLGhtlRvvMJvX0lIa8ZMgTOFEPG9O7FNARxyG/wjKoFqDf
6HAqvP8b5+97UQizFkjaTx3I0k1vNpP5ysaUSoV2gPhaemhqeRxdJ5NHbmbGyRfX
M+TlL+uCMUVmKfVeL/do1eHUjeB01BMtJgntGhFGUyB+Gvhr4HVSdj9kZu0x78vF
PxSrM3mm9+il9Mu4MNtFi5fhjDZolnHE+ebRRK1I7N4Q8/1KP3IdqpZsKIkqvf1t
AmdpDmxoyQj9jVGHf53eIgQsHI+mSLtr5U4T9nJORGSGSyY1MpsNTwGax67xensD
wyz8DFD3842c2dfuA+o67koHB4Z0kWifIvf/WUamCH8X69QPD7AmMWLFAWylvMun
ze6QNbY9wrL06DUcqc9TFXYTT1ExoqxBMEGzXA67BRh0IENVbG+j3DpVytjXG1CH
6IRRV7tEFo+SOeDrM1h6PwYbqkB4/FkKjuIl1BqPziXEP2KyF7GagfPWtMxHL4uj
K1xvNSvjKVB2kljjLM+9W5YerxcrveluLnKHvJ+Y/kVvtzbpwZTYjbiFfPuavfZs
7MHkgG6qK4HvlgKAe/h1+8utrYJSkdywR+zJIlJK48lB/ZMqSmJNTjxwwbwGvI7O
b3sr+Wj7hpxH7R+Dh5pD/v/iO5mag+HiuLFPcV7SgBoCyzp9yEFZZPEWdJ6N8Yaf
GjGyFH6AJqYgw4VVdfi63K3vKt7n/5uKCOToS03AuCX4pKUKKzBFLBtJhSrM+d7b
qyPK3Vplwxq8EaX1Thtqa3M6bsqWGEIB/dDCB7GR94BjvYrNNUzMLsHHeOwXwNVf
UXI42KSfr2ARkkfjuNGt88meRIwVOeErYMkRWo4Lgq4+VotjFMGVbu7G6Im+XJl5
S/6Lh7YOJSgRzJe8vnTAleKPJCLPoLSaNGdivexngBZx1tkJtukQBAxpJaknAR3d
WccyvA5G43V0jrRVK12KbLPZW2eGcAaX/t0jXQ0QZq3ElEJY35N0ZUkDiQdjmqu1
Ii4rquaSW+jnyE5kcGgsYAPCZIE1FRYr1aQTEsVb1ZvCO1X133e3htR0qq7JsPHZ
Vy5rLDDoecjzILbGl1ef6ikLkgm9uxZPxvlYQVdnKTpOu/f7/KC0sS+7L/kgrAHQ
B2C9BweQl4btzAu8dAeFcvczp7tZT0XHGSBxa97otkPg+eLoV5nAJmN5JUiDdLDP
1gZAp02m8Tv33WaDKQAGwcZVIAIbYcQXg4gKeVc5BL9T+4FIgmr5S6iJ51uktjx7
Yk5rE7xKqCJ96kSIqcjs2UAiqHKaKGeTN4eIraxhL6F/2Fqzpx8CLeNgyDSUXZEO
/KhVhRPrcNWlvs3brkTyyNMHr9Q2yxdwIbGQPNl7dIcU16NBYu1boD+b0r6HNGzG
O5x/OgFhtAGO2FCNbjgMkdSEiEpFFbJH+EBhJiFGq4wt6P+P+txFnY3OriLSAFDu
Webm7pZgLmU56U/z2wzKTzFt3z68nPwo0pnf4Q6lYV+l2pyK0HrrG7lSola9hZBR
+MG3dbBe1+uTLQH2RH4BYpupjGrYQyOlIiyU3nOAZxeiUb78TtmJyNdrJtxvNJRN
2PksWoS+p7OHwwI5vIPmHIPXXexxYfM89y76pTCi4BwaRAD5Q/GNA/hdRFPuOIc3
Wd3I3q7wtQGgy/zTAtei6yZ3t81WUNM8qa2O417ACaf00Mkb/VK2LTTTyR3qJ1x7
4FhecqclA+d4rT9+Px3UY3D45SNgeneAsdbS0pis2vFLqLE85/efr7TFrQtMToqT
t5mQFVJTd0jXDUHh6aHOEQYETw/5Gi6XgdBeFoZ67OxxyeHE9Fnhg50KtVTTsp20
2XmaXgKFoNZiIsaPdywV/WtiYk5tSBP6NVwZZ1cWwDLOya1hnwJ4jB9K9mjXCOvM
R5Q/olwk2J1iguLM8jj19wCb1s4x+dJuoZLYA179+zNdDEUgfFSAPNGlxrmJM+7l
ZCIo6/VIXOFqgtlekRzzh1bMCWNa/TtYnDmQSeSEvvao95exJSV6j61IOm2GStRi
4KsJ8Yvp1dllWuJ7JCXcDLeW4EOuI+r81h7P1/qcOSZtBhS0skRaYxGBMrNA5qNg
eurPa99vU2bcgUQuv6y7pd0xz/qvX4D4Z4VGsHI8gQa9vn+5GTGR/cee5OAz5/5y
ExyFeG5KkxqYAEUKh62URcs5kKDQ7GpuLifi6dVXDGZW6gMlHTI7X6eDf5ApTTT8
G1ovXZeQFoc9zUh6lY1eI19n1ORq7t7xux3aH1p66cB5zOe22ZEughOeVmOhgNSX
6VRsf6Fs9ZvSKNjl2iFP15qUOPWsBqbq2F11GxtshT6e6M9CFXuFIdOfqZtV4o8W
G0Gu0zo8+m2ty5HN9ATIlwSzFQjZsXt9yBtCNNlsgYTGVA8Ko5lLK4buPwOF29v0
Re3ofrLTCcGO2hi6ZI3pAzfRqw4GUAgd48NqZpTNpr7z9O1S7EEOZ53qvvfMbh89
13/7mixhPDiteMsefiW+1ctyWu+Yqu38KouFoyXKD0EfKfPGqjYdzCnlHlz10Nq4
xWvhxcIvnapykuljQK0miexpEsQBp/U49LlshgmktzEYRq3yTs4FWzTBhfvYYn35
1T3qVKrjMOS8dm5qhFngIe/FivORr1ELY4hj41ydtTG7XWE6sx90j0QFRUk7UooK
5kjvIU0JW3FGMNaCqmiF6b2Jb1JLi9Ag9xuV8dheZxZulIUCOLCHPs3hYnNgWEIf
naJj3xFb20o3SqMvnKPmE5jYD9GmPHbprFkZk97GS0cT25JHyFQU4O5Ucs+H2ahQ
Gr/sUfAgA6KeD5fGFqZ109Gj4xILoR3czgsWiyc+fxWu5etpNtgxmFeWQy5KkaPm
XyGcx+jNJqVj9oPg+MaF/R5Ye0UnYXuYp6OAABg5BTS0Lp6JQS6aC4QmpWEfmEPU
Hy21UkfRHV4vqEEW/s4ZbycWkoH/0v5pBZvbqZ1FDstFvZAU4LZx0/yVuUN+hina
euLhn5e0lwkc8kFH3BxXlLonHN3Z0EosdImYHeUmGneKmyqj+pJ92pKMfdVF5izr
uApGrwqXofaAHfiENOKzgxzhigLnQcc7wQqyPk8Zq+7x33xFvw/S89QtBNYVsZSe
y8Aq0f74s1UgdICmyjcCkYb3F/p8Z4S3WURLtcnlVguVbLZGzwG3TqpaIro83W4f
6k12k2At4LLHG7bdk57JuvGLm5l+v6PCfWtK0xtxcEE1c2zRqEoT2DxDhqDOHtYl
UApH+fuBBBz36YhQntTR0Zs91uRqzY65BqvWo0rbkuMci38Ne8+UJ+i88pxN1MjW
T5XxZA9mcPd1E1pqOVLMCNkt3xvnvLWMgXW3PdO3O/3x1NQ7QAvM6zJ/qtnOOJ/s
y6lvmd6uYL7qMe8VRZLE9lVJwyuDgyOvJapKe5V3106NUYK10icb9XQdJWmszge0
Dt11al3DYYkr8lHSBlTNY/3SV+7ulZfy08jQq/Hn9btEZWgIp4DmC4QGOS2PGM5n
7qT5ZqaZGf6HU+yGp/zN3rkoE9EYtGMuY237eDfy3HCHj86bYfYKlNbWUW9dfgmY
w5enh9vvFWkEqVVyNDOq+bKliqA/MC1+R0tAT+bXtdc02vmArYfP+52wUQcEEjgj
0wAZSNGc4J3OKEzVarZZro+wwy1ppiZun2VkSADCCZ4yqMENITLip0DAcD46I7h0
IO2hNJwna2qxP9F0MmRCtvy4U5thIq0hLrThRFj/xaad0GsSGbpcI9W1YdHlJ+HF
cpluU8M7sGZWGnE5xSiijBkzgegCbNyMJ4lIRC8sCP9MlaKBEzRE+an4ljMfrm6p
yIjg/B76V85iz2jHwYsgOOIwb3mTZ3DrJZrZoeI2CGjx3tywpu2DxQ2jVS+RKbN/
1zxwjYJ3v5nPFMr6bRTMhsGuXbasdMrgQPndGEzMBgXoXpELdIBQTB7dRZVdaL2X
HmqG9wPDA5l9/JFVe8lMhBd4C//EVjEE+I015anlgNiuNrbOTJ/oFVhJvy9MtQSY
I4XPFUiYOXoGrqEjKpRJKcO20aQmlvq0MvHyGmkyh8lPfcEsQ9lvkxSkbiT9zVJA
EKHtwl/+giV7whKYWyaXn6eXipoF9lTBysaP1TtiTpVLdmnXKrv/AG71ojeOH+e6
2jLTR5bBD6jtYymD9CiEn5eLLSSFJISetXt+uXX+Ln88N1jSV38toFJmiO/RTgnZ
kCnWXBuIbfQ4D8+1E9z5Tndj4AeKPj8yJTrcjmFLixQ0Y72tFcPsc89bRMV3+XxC
6ZDHZTBm5D92TkeEQx5vqhzoX0z0mc5UlILSz/bzPfAky3XYofSuy0ufxj4HHAUA
Iz5h8QFrSxrDx2voQlZuOCHRt1x8Utg/KZQ8aPLjjnap6bOJfZRL2HOpxiEk3q1I
umVj80HY8aEiV5mPli9b6JxalqLbyWwGI8BDdNcG24kequoojgCub5Fwd/XoN4+T
BfWi0ak3w2D/cXR0aB2qLlRt3k0/9PXT4Lw1YBtW1KMvwZJOhTi3xciv1obHfMBK
3YrA4HZiaglTC8KHB8qCcyB942PopcB3GW2BO11v7dpk5EOLGOWXaZaOYSO7bE/v
p1wQQ+iTj2s14dWOfzDrO3EvFW8l1iGrVTH2I9CTJdbsltjaI64pEMr2YSlpeX8C
VS84EQPEC4xty3Q7WdwuzJe7wrZMqvQ5hKuoVkGd7QQaoindZgfjb1M1CQMM3VPa
imBzP7RfiuOBZgn2bvhuGoKPhK1wn/NXzEFmaXcH5rCNRomXYSRQqYO0NCCgbK6y
i85OZUZNFt30vO9Uz5LbuoEx3oTHb7/4gJg3/JYHE5VYEmih9sjNDuIImHjRUHYN
M1n24mEp4OcynkxMJu7u+CluIs/Jy0yGBaIZZesj6b7jSmt0G8DjW5kPPZBvtCbo
9auHacp1NjpYIzGLL4NKLU39uShcDhzg7kgeHR/hXOsQqAo4zKGeFxzsC8l3P5Ph
K0AeIh2npzjyMcfj9WKrxpmsKrur0yI32I5cQnBFfAroHOTf/JFWrIrz1uH9aQlD
uQt0gW+vEO8qOgbuw94dwQglCJDxVWN94iBqgXIfqgXVvelH6U5eBEq1kIJBTfsE
zBf4bPO3y3xvynnKyey5uy2/7w/MEGHPosw+DBN5j4xxiRc/Uix2qPE7Uzp20zvd
iS9R5cBDi1XytdRl9aNDrEoYoipGbkdnA4nljVySLBDJXQfaJfn4Kpmr0MuIdevN
Ao3N9CnjqAbiYJiTw3DkVwMbRYleT+6FspI4qRTR/b/ATxceGPoQDKVT1uEgr085
Lx+cS9RpSn7yQvAI0LJWXVPQDxvIabr+nxN7k+JGKav3fB4IQYa2AS5fh8DuktUM
hqTM4l5T9qbzAsckK8T/29YREGONIS61lXrtnBLLjaY1q2RBjxFdB7IVv9IvQbxA
tqerSJAWXw/NmASM2tcR1NKiWXvME8VEqDbEe44kdR/0G62xK2bEbCkMTjMoFoUj
q6+krXE0/mNJU6o16vr3mOfzaGCfSTNKgpho/t6yKpm15Yws/wsWMEJ5KpCZy38b
K2QwSu30Q8lvzM9u8IyyYJkossEFidqShMJ36IHMWhXF9wGSHZ5ppyJrvtTp9WCx
gnOXOK0th2/EbxdeUglrXdg8f253RniyD0U9ChVKcV4Ve14upuAOJxjQEFmmAlJS
MYWxRKeMRnCodaiJb4nkLup+QyY0Vw8sUZxEdxeB0JrDBeSYUlJNdHLpXYQ81iOC
Rfosmxvfh6kiWUFlhzdar5QNxrHzPrn//JeMhTOkwchr2GtWV01nEmnRwQDUjR1/
yrElzwFmNwrbLsF72/pG6VRZtIcDCw9ewGHe+TZpmipdfCgq0w9OiYXRJA3TYsw0
yG313VoL6dmYXbEM6tHQ9CCytVOEXUFkC6vGb4cGCsvCIKows7zpFj+hSrMc0mJo
hMszssDE2P5aVZwAMoq0iE0Lme6Lmk94hvx+6aE6YiUn1YiO+0wR9wZmOm5fBfbb
UJXl3aO6Zh8Vn7faViL9qNUxBqThJJIKutM0u98hyIzuMiNOSpJCHgd40Q719nge
8QR1/xiTbVG3ce8ldmjWSmfKZ0Uq1SO/Znj9Pk9T2PyWSvtguxLfHRy56VmBm16B
+dRfGjtfsthKK6uqrGSJM2XuLteilPz6bLzF1pz5KyHHlzc/dLrkfVspH2HgrVq2
ueX+N2OtUAC/UZD1IqhVD2mk3ED/umKyHcchvPKEZQp/y7J0gK7u3zeJyOWgUjaB
hV9lzVQH6IMHY9YtauQQyDD0XonMuZZyMHqKj2krW6TSGOubnVsc8wwUwAjXFKft
NeTu+utzjPf716bBRALH/XHOEoYihWp5GvmFHBSJcmGhkdDtfej/UUvqr5TbeNy2
guXqcJo5MK4RMzb1nHr5FTfzVxrqQI6AyeILYcXKUD08cJ86AWqGXW1cauqenhG9
o1e16v23uJU6CRM+aa3Itd9301o44GMr1hJdS4emTiTAnXLpYROSJxYcD9tCXj5l
xXe7ahZcIf1Qlloq1ulsbAWdvzh4FS2r0HnWAZI1mUgqLSH5ykXDzmI0uVNYd9TW
jutbOJ3XzEiIL203bkP9pNQnTQn0m6OyJGs36HblhBSwd2vWq3/1xn6PKuswtIty
CZe2l3MbDD12I1QuiOP/9P2N6mPOvNOaTiIwCoJQR8RiwHdBJ0p0qsLjbXKbhNtG
RCtDj80844qlEG76MqvalwhhDyIIi/mHnRN0aRia4fgdmpHwgzAi227UZU42RKkw
Bzn+3bTdGaPfE6VOIzUxoWato1iszChMErw90mMn6R6XzuLq1aaR3h70KEeWFWgb
Ep37ye9bWeBnTuYPZPpie+oI8z4z4bpq5mkhb1WoVudNDWbGcdCLYRXIG+UVIkbF
Nfin6dp7mGg/XNNEo+pFK7HhV5wKUj1BCwC28si2R7+NDRBTmqNeRbdE8UUZ4/9O
yrlfM8ipKxIi4fp7gOfmUQ0fYzTiCVk3Sx6WBXta4dUjJo4xPlgTKXvNs4bql2nV
rTucvU2IfG9qk471wwQNiBkwTeAYd4BDLttoYy4Qlgkn5bEMOjdfeQ6CmRK1KAJ5
T64MZTNCBuJejtVUekWbhyV6F2/gAn1OngM4W34lBP0+2rpLamoW7ZGxy6K6v2aj
1PKomUiW6zQ4OAj0cWakHcMUaWKg/gficT06M7GFjhMtLseQPPtYX1miAZCW/wve
uH6H1ovXYLPBZpzw49RpfElLlO1q1SMHFlh+P2UkOelNferrerCEvLkZbt/JSGtx
q1XjzuWDZ8Cy+AxNT1MLsCKnWoTiEo4IMxubIOuSmPYi1MqxZFIFO91f8cSgTg6R
w7+69b8osD1nuywc4j9dCFcMeueStCT1EeQqSKguxlAgf/U3h6KJ7UwQ6FG4IkjI
enB/gUx7uombrHeylvgVhJPkfedU11KfaRAUj36/c4TboF8zViLFrUjLOaMBDECc
6xPIWSJwvJ77TR3qeUIYY7FbUW7MHvtII+gw2P7nkbbfM4cI1ku0RA5RED38JesO
DPO/PYljOTdKQWFEpPtPyuM0JbbjiLsddbmGMutyFsThiR4nYR+sUUVaIWKGh6/2
yDtbgfAcHq4UWkHw+TWryhD9MSoIH2d75gxow8BG6IFFycUM+aMUXSRn/tOYJxgd
k1VdezkBrD3jo0RTi90sp6GZu+xC+HrLgLdQl2Iro9v0oJqMLNiYqCaF6RfR6+nW
tMTNfeJddhs1RKl6LdNcvtzbedhQCcPkKx7ArsOwMipwPmllo00JLpAatvLPLC++
xeuicW41zdyT0g2HuwuGlFIvOpvZ3MKQC60NHfPnwLTyJHdCmv35GrZweZJKUIj2
WACknGavdDcoSxWDh0EDhBWKWAhVllL+CKJi5eHJ3NZw71q7mtYW1+KIYHiDRR/W
rgzdh8ZW8y/gYTIwU2R9pZiqnxNtivvpzNIwX2jv8kcyFimNWyiGI8iXZ5h4srIZ
TGlDgRZir5Z4eaRzdCJmYgVKdARA7RDMeVXRa6dQAe6P8SXs+xPO7M/mhF107MIj
5mul2aUeuEMoTI1RAJ6x47VzXwCLTnwWVxkn8Av6yXH7p4Mb3OufjRQariyGBHjG
KvLJ70/NdZ8Khl9WpexA63A22nphqz1Bzp4IBEI39q593TU8kZoCyp57P7sDcjIt
yZgvzv+sa/lcZQuSBs9WEXVZqjBn5DkK7KTl8Goo0hZA9dL7doVvpSakaum6MPOk
1Ry9IA6W0upbWejkhC1qxbDv68uBm1odERGC/qGqGCZZx2C/1QqA0ZSRCc7sbdnA
SRvaNOpU2MR7lcBG5gy4//H3vFpWNZf71NYf0X/GltI+cL9L06I1hxFGEZ/iU9BV
Hj+oAWJO3HDzwb6la6aidWjxMFOagnLO8VVDW3FlGfJ6eKEICPcPauyajV/arX8Z
elA8VMYhJnQUpo2i0fmihg31fRYJ7DUzxdyvu7letbzHi6bp4ClKR7cYOK4La8wQ
/jelWYXVthlL0UwsOF1RhiM5oaCo2kgPpcmYxiJ74sBWcXZq/bV/HL8tuwAYplT5
2lrb88I7zDIjnza/RU4G9wdpidSAJ73zxYyqQTQRZeWykaItvbYZ46F5X81wx4ch
qawh8jkP6Xsxi3JQ93/Fvx3/F8w/PF6sObVJXwVWkCCJnVtF09F3Lk2MSkMWtWDL
HpVjiOd/P03gNjF0XqcJWGjupx/1lou6bU3/UfuVBDeQONOW0Q9pemRi63nUTlJk
mO39Ro3P5g3fdIhlYDv9OIFmwv4ImkQW6dF7s1/IRGAuxhKXbiWpb9XTUTaruxSO
oE09E+3/Io9CwhWj03FPqC5BhODVO8pp6ucNNs7yo6t5oakoxaqGjgyzRwndKD/x
uU6fWMK5O24Yk1tQ40nzvx5iuzN2fZS3YlfolYGBLfPYbERunP2URstMWbkWLtI1
u+ErgUWX+N5UzUiFJWd2plmQsET6qGYBkAmFWwh+HkupvCtZ/cFY8vaVfGX7xedH
1/QuCytuwrkteLI3btMehx0PXzISGCfcHoYc9RYsfRhsZSdoCzcDkQD1y9KIrrGF
6wgSUksHvAk39WRwx7z0eVjR1KiOH+qEKb9C33CXi3dJonnl5p5DTTXDbH7JC7Ss
T9Ar/f6KlQw0jaPM3bx74LblR7b07yT3iIiqnqAnE7f5HdHdr8FEKMNG95aJGxyH
ZqyGrzM2FbuGP4mDGMdk8+TbsHG2JD5yqRzauOe7EFAXyWW2qcQE66MLOzAqA3UM
rRpRL4p6lU+9FrEj2d8qXP2g01vDbGZGa3fvRswzh+iQp0DRWFEE8my36fjOqd6Z
88LjhJhDyqAQd8X1Oa1K1+d3t82HAa0YQt0bGBBLssZCkVbPM3MG8W5DCGlCDYNC
inwc701aBbA9tphX3e9lFNb+bUy95AHR/2A0pZ5oWC5k6u4F08h/zMbVkmcYZBdi
pNYhxjzKJZsN8QuVU8CkWUMcvZI/TK541DiRI9Qa2rTtV4R7hv2mscmB/N4EPH88
ymGEX3E2FNIPm74kaC/1lrNFbvkWl7hyd4ZZ1mHuj9Uk8NO6FrJs/M0LHKa+CE3u
HFo+hhB2RtjGwCiM7GstU6VKH5R4oYQ5drydIRCgDx13H9J9XC3n2r0mkWE25JsG
D95ZDErJCgibZAJomN29Sp/4AmcPAf60XDqEgEKEmfdgZVBHezszi5uVXS+MDY+/
OhPftqdmAooV2OUVcBQWMijjYsbNJVbx3CsVkziN6RhEYIYmM1GCobmS9JqEGXHN
gXlw5lDlmecUg18/u9Hr5pCNQE7GP386QjZzLGnhWZYiKqdgfX42NA6KPbQzjXlh
8gWjSeAONtMWriIsZZ347/Vm+d728ku/PEMrNM1RlaA2Nx1vRMxx2UbCcjgFteQz
BCTDieFSF1ujvmvLce+eYvuEQBzOkd/XsBrKn1s7+bw+j8Kq85emeuglaGZVa6eN
a9N6GZvkSeMCvF1KybqiOs5Xf3DPVNLqBJJPMZDGmCbthi3NXaO14H1XCIVk18Me
KElgSK2imXwiH08qvrIvmdjMpVOBx8lqqHluaLWnxV1rTvom1dXBpt9gKcZppht6
FGwbwaqW8kwa17Ynx2Lm5ubLaebeyiUT8TFpUWLY+MeDsEKauM4ZeapmKWWYbIIK
TiwZuX9Sl9lHIY6AVGENnEFCG+brbxtYQBKHvBVvvRMXJE5od/gvomoEtwCDA2CG
CeyhYCerPQ1ZEs/DNnostfDoZnT343YuN/6RNJZ9qD3WguX+lkw+WyhRUAyHx/JN
x3J12hk7+iE/ON4ugxpUEyjK2DJfmEQi0vdm8IVNkF3lzv5ra2aBNjXig1A0PvxY
PiVOol9MmenraTZOsfwyoIi3XirAAmObQNKGaTS3MeDJDo8MMHM7ba5DLlnjEVV7
bnSmI5ByfVEsw0TA0xH/e5UoBD9F1+tANvjn/tG6dkptP19bdtRxvhm2MK4fSnXu
/qfZ5+dI7Yijg1gzxqh+29cEarYuVW7drrIA+8CZUSK6C+mb6GrYJhBl120DvNvr
3xaOjhPeJGcaXswuQIEQ2qyqHNq67qqcsnD7wDs/SxvJ7OQSyhazEc1/001Ma1CB
ro/SOp+uWVCpKSvPrR66z1CNYVr0OkEq241YwQ/CuDFRVJQH3r3kzKqTEcktr6R7
pXuTfT/ZCTA+l+t649Qwp+7Qnyu4RwpPACpnu5ac6Y1wcQHgdICmYdAYODO53FrU
G85wL7dO3oiD9RdYwy6fXRnN3JsMcS2pZS1tCY/qVTGCJ/Jn7JKB6BIwfpyfRq7Z
OKi/ebnVgNrmj7TE/JP46xfQCASuyNfBnBG1v4QiMQ0Bfm9Sg8911pKiKcfmiCDy
rRIeWXF0hAgtE/N3Ynvygt0jQLU8Dvc2IKVNqcAe3kKNjWne++b286uyzc73oYZE
B7SOE1P1ZIJ5c5c2P360uE5c9raAgtqg4Jm74JB64oeSYXOxuUvOAOK51PDm8QyY
/KlIAa7Do9ym1dckJEKxs2FkUYi+KHKvqw44HTE23zWno8Ngn9U2C/lYRc6vvGHk
VjoAjkzv4IF5oYxW4DHRPKrtEpF3tTcP6D6HtvZkwMci2f9i5lBuPnAtd7snyrZB
36HecICng5RprLIhiSLPBDKIfvu2Fjo2WTCD5//DxR8UTCK1E9zUSnfDV1kvDFCQ
t2Hogrv0DNTURU4oNVJNONPJYCSTL2AoXqCUkcJd+zvvFXDIwnyjSrxxzS6zVM5g
EgNOs33ky7r8gDt5qk/+ZA5lR+LMnDHuXCqHX246dV4w7fb62DAhfrKtF1f/+/MO
d8MU6Br7Rvf5/bnsXM65GEtDyO5WBzwCQanYwOyGluo02ccjzte8ZGJoNU1HK1wc
hPrHm4NpcF0VpGtS9atuUxBmyMOcV+WHxZqLJeVak2oaWdA3ciJWXwp7cFNHVCI/
i2uE0FnqGuTpZS+DOEXMcKVQOHYoG1zsM6loko25+ZZuYQ3ue6vz9CGJ7Hd3K/yE
jrGOGhJv+Y4u2ej2An9EwoCGfKl+bo+HqkvpQqup0ILTUIHxkjlIF0+1vglMUwvk
dZJqP7SSLsEsTViAME8kjX35uIGuVObXzH0Kj73Ew2rt5VxZFT267UpQZ/tSpeyJ
zGzqgkODthxEbya8/a3WWtU5S/CxIwAmCQx/2k/dvLaQSNK65B3rSqfLlmX2zxMH
cXr3jnmmiwp+hca5N+T1cb3BE+c/9LrfHzlxgUiKNz1QULLKoI1LbyCJpFXvoO8a
mRIqKI2RJhXKBV9IaVjqE3/u3dlSEVeGnstXr09qncx6/FJ0hoe0Xng1tX8k8sCJ
IpAhkBjmBd8AJjOLw2tTuhuvXjNIIlwVEVrzISvHLtC2pMdPc+BEldVcpl7otgPg
XSDjOO72t376Xq5uipEqguY8X5nh7DgLa+buJrNMBLN52S/BAfv+BOvw7nTzQb4o
v4H2qh20atVF3/gy1PhrtafuMyAJqoinW3zf0mn73twr3I2+F6kgcZOVghAqCDKM
MxUBKc5TLCOX06N10TBFwy0a1YkFcBnEXxhuyQmT960/S85YsNFSPQKFMBtJPO2X
/5ISGAbpmcrcQwUoRwwSPCpd7Uli3EJCCvTdWGfvDUrC2m2AlExm2QJj6cPqoO7k
aPFqgZwvVG87Z2SfQ2rs4NLvcVcEKswjW0iGwTs1vyFxpDMdxizGzP7H+Lp3xrlg
KmUJHA3gPsmexDJwR1Rz1Rxj3KyUhoXYgwC/heF9o56ztFL+ehQGlINuq1+ShIcx
nrAfxDnAH39veD5x5TkY7RtYlU0kXQ/+DTaGd3vQN+bDPjeluosAT0wDjayJ7FWJ
EA/Jp+tgYGX+mrO8LumHoY+UNc0llHLpGd401fv6nmJ96Nu0nvFV4Za9QPHrR9D2
9iAO4lQ/sUnF4iVGU/PzMjjabfq5jDFpUfAASQMxCJjWDxKKWgwq8raYKrIUQI7h
cyWpkj/LjHsxOGEey9ZIyNHwvZF4JTLofOz5OjGp/+m8exJo/xNUlPXjLeDwnDDI
2e99SeJ+n6bnTxk5FWOUAtvYR8bCCOP1EFw1f5v33nciq3wsZ7IeBBnCLGiTxsNy
cuYsJ4YAdpCw8rzMTP2oGHVnLApWRQT9u6klKqwzDdNsdTn7JumAv1W7OK13fYuo
t4fOplHRG+CBskeGZfxKwUDL559XI8rLA8EsC/F7/P8bXfHJQSbcQqIC+apOObts
3lBE42Z/GtfxyZNDBTldATTq4mKTXXjctUe/p0zyBeyBGREglDNiWoDtDBQ0FgQ2
Mvdtjkrhk9P1WbUV45c9aL0QsHOV5Ee9Og1ujKwO9V231nTWtcO/SzodrjJH7xE2
CAC5RIAi4xwNFL+P/sJqYfDKmrI2PhvYsiLy15djTotNACt7/ZwiAPG6TDo62LBQ
qEij0ZQGyPWgjhIl1hU9/s16ukDWsbn6NtyG2KSVBT71hT+Rql7TXE6Yy+N2GZ4S
ZblCOFRP6s230+VdROpnJaVB5Gaglu+XAHpWkFDliK0avTni3G3tCsZ++VvLWHL9
KUpG80LBd7lvqaV7TFSTzbUMpauIVsgn+m+ft9YKkiHyp00WLly+aMzOVrxpabbL
e1Nah6hvAmZtNYDkFAHALXofeScG+VGMUo/2SBXd0FERqTALcLYeIp14ckHPyS0x
RIO2gOo5BoKggwmTv8+5i44SjpeKuGjHEx4mtof3F/oA5WPQ/5ndH00cU+A4gs2X
KwUE9IHJaKvxTYltly1Ce8FaYBgFgL3Z5VK+KMOHscE2mIT2j6q216jLuKZ/oyVL
NniUuyd0LRXRgAVKhEJFEvpAH+SFlgQN9Dx4qThc9P2/kue0S6jvpoa/DwJsjjSz
2kIkEVhlidh0csKbzcsLqlAilARC0MhIi9rLu278YQ0+K5miRtV8p7Qqz4CGgcAy
xdxlG7RZi3dc2M2/rhQyxbKcyCAeUKGV6DgbLIDZNg4IGCDjc5fiY5m7hHgcD/Gw
zcB3WHH0ipuSCsjqbYrNJXBCJWdqPxAMWXESlD+NeCaSzoKo5vPqY8Swxa33SWNl
9AHlt9GuL/EH/RYCcOZjdrBLYopKVluL/gQne+S8j1qKDbtXO2MDkExLXih+JpoA
4b9fdKXdc+S8LNEBcB8doRMz2Z5YJ3iyKqwyNe8WybzVYVAn4sCzLrR4nQphby3Z
DhFTLNfI7ull8Mw2FmDT+IQAitKAFgojpEWTHHnsVTrWkWMfOB8pmom+b9CJAW2o
5h81DELBlmJZmjHCCnUIHl+y6fB0fTzmuldvB5gyWrZi2UHadxazWTkXEERpxQTH
NDDvXd9bFWJKAYynfV+3/iIZo5et2LgKL0l+Q6y0izDT6bsFmf1ETkGBoo+yNgP1
OIr8UTqC/hZj4EIgF4K9aS0wHh2DSHAJ5H+f1fcQ7RSIjD2jZwagxMP2Ok2FwJaM
6aPfQHQ8Eq8spXuVHDo3cKn6kxat0Tjxm2/UTIIZJkoIryoG+4aTcSs/AM8FFiIU
qlrLjWTEh7hvd5KrtNkZ/AOqGBqANUW05tCM0rpQFcyFHgOrNe9tg+KKJPrJCzuI
EZO3NS8sRiCuTE1BcvNQEQnQSWvtduFMD/uvQGNZmQuCCViHMNLuoacJYDFNXFv/
t+wpPLGyrL9sp8jHAQjiidiS5U/k69W3OS9XlcTVUP0rR9KPiMn3PXm5aEGiH3hL
BRg1rgiAIXEdwGJfhcUpWuelM+cv2y3wLh2fkXlPfmqZX3kFD3C7JLN2Qa6QnkAf
8VWKPqS0vO38bUwfYvuogPcTS/WdzuQGSm3exmUHfZZvtxJDKgEqfY8zmNY+oxvK
J6yEmtKt/MQ+ePgQaIpUesQ31J+IgBIEpDZ4b0EcB1ZKmxh9P7qD8eVc8/BpRO4F
xw2jmqA2MhUxWv195JcY26Hw8yse4Ir6S/Xwl00J6hL+USOLbA/+B6CCnfCboPOa
R434U/zHxYOCmAsHqXM/1w56lOT8qLBct0SZuCOPpIwjrlMdkt5gCY32uAQjaTd2
GHQcDUCAA+kSXfc/snaiENfuYZMuGXSkqH87x44uW+2Krx8dI/GtsNfIIjOmkPaW
VMzAmrvsCstI27PeOLmEroqfiKfqOKzUGeLOm/G81st/B4cjQ+YdJWRpTH458+Sv
Sx2j/A0mXWxKejyhruRmOETNRV3VwE3rfS/xyQe2xPkYDDBZLMcTOar8u8VLaZ1c
xLWnwkWjOf0+fIrPnjsStBu9k7ULL5LgtkObAEj9idQUjyYFVnBjm8jyEsDBGxw3
xXZVlD47YJFgg8ndCE/YcSOMm3n3Sx6voD9hD81lXQ8y3I6CvENEAT4f1IlSbo+l
iQfe1Qc4AlikKfn5+nikAkRXDlDUOk2KTjHfZGf4e8W4F5WQ88neV9OVXjyqniJo
G+K7mztWSD+JZEsaVEZzHWR64zrkVwqB//rDkyoab4RCq+TTz0n+RrW/I+QUMs2Z
jD3N/uqt0ZfNRg4y5FUkVH78KoApDlUBjpo3UHB/pQZJGEBbXPhgGXIADoY+aJqd
uv61gKL0H4b5vc8hezk8pt20UaJQqUqV4c0lstlm1FPwZlD1HRF9QM8llHFMGh15
ZXTSdqfEbAloJCso/BSEcKKIKTdP73i8P92zNTdCsWSYqAMvzWws7UVZ5/hfk9bW
qEfbGstC/Bzsn+dTX8KcL+zwDwSk17Y2RMQqlfRiFMXaWKZmGo+S63S0JNfr4HaX
cAOt4cRH7hKTXFNTn+88jZSd9g8DEzS2mFsMi9yvVuahiWsh2Wb0AHyYmTNqYa7J
L5SApMV5DUjmmOlUHVDPBiI3PSJuSvBvfWw3eGsO+HWBOElidsnZnwZ7lZ4IPXQ5
+1TYN10dq/z7T7zFp5zZSRsnhlbdx6DhI99auAZMQsS60Tqf2zilnQ0efAPrXE79
FyuVNch5QKZY04mKJtK9ZmDjpn2473U7iPhvRJe5kMvPt7cs3wSB9/Me//ff29+7
YC2MuuaEjXTJCm3gAZHlw/gwlYHB5WK3Y8eZLxzo9piQx+M0rTQ8ONEa8eqX+a6h
iQxhN9oTpaf5TVj62j4gwDwsfLxCQNMupaNj/NzmnQ11IxNoNUB4hhwOC3NNZ6vj
kPceRdpnNJ5PTSZCg6MZtRBKWETzU0M9KGHIMDsm00FRax2OsTf3wFR3bKgeQILy
+o5wBcmQMoX44AIbkWXo2TpVuArEwpZxLzv3oyHwdZG8B7jkwM6IvAARfr2kjoiu
raZt1L9RN4TE0KibmUyXIepEdWYBCaLL7IBqyJ5nuwhXj2aSXtOKiCB+277u8php
cxMintiQXP8n435LY+CyOTE+h5TTmAuZ3YHk23AEfoTEZDfpgNsu5jlP4BqvU/ew
gz47bu52eq+YJ2bax2clZJELt90fYTYyXQhDzB+to7Eu7XgDPZtaMJYHTuI5LXue
JsqWC9KUP/fpi8vjTJoavRMEe08t1V7tYfoQ7QZQIhBuLBpKIZayVUJYCraBW7oh
liLdscHBUaTsZreyPUvxJansZDU0+p3Kf+VMoTtiB5FETl875eIBxxB6kJKC0KzV
YXzcz7931tmCgc0Df//u7l7L2tgtsE00ehHXEOMCdgC0AqXuQ8WWUkeuNmS5skta
SzT6JgZUIhcrOwyEXM6nEkxfVlXTSw9j1cEaQ2fweMKXMYzyCfVbHB31UY65zKgk
857f7PpS3tjxKY6f4vgFEHk8/l11oRCunuVIU3xi1b1eu/pbfWNqRc11yXIUXLBJ
u0oG7YGVE0JEJVBlZtGXmXETO5sjjd3iI/UKDdPjeLPnRM/ol/7fMpg4BZoIAkkw
M9EuxxM2l5SbwpM4bHYzv306y86m2rS+AssWnuxcaR3fiQ8fsvqLwSlNvV8MSu3V
LBkYuSB8el52qIiw8Mc1mDmjDkc3gU47o2Bb2f2sjBUSalIST3iocumc1BoScDO3
EdmI8RmcZSTMSj5NboSaW+TsoczxdWPVINXM2wLRCpjxEQQtJ2wbcTyrnBI60nML
h0Ms+3LGs/HvZvwOfQZ34v6z3W0KZsJH0itPwkejmmWDg0eCTh1vkW3x2u1Lk7lH
KCOgL+Y9/caZS/Lt2tTP/OY80aXcct3v0c/8VRUsK75rFMA+Z4Vj2YVmdg6/cmVa
u4b7xEj35eqYVqWswPoN88tP+vXEoY2BeoOVA5T1SiuPQV30C4hseqyEUDKipsBc
vo7aFWeq5OkF1hwj7Z+2IWjG50IrpTiit17Jqn0POJDR4wNKPjv7VXWwFtoy/2gT
aj1fn2WLeneRdN3tVbm8y7UEYeD2PVq4nc5a3ZwQsdPYJAV7kWN1A/Icw3CkAZaL
bnQcfR3OsVF2i3IxwXDRqAQ+UC1OibTh8Jxs4KrKPv6rsTHBrrHxktlVe+ESK/wW
czN3w4YR4E42sTrhV0ll0WuVkLs/6MGpZDNnWmap85MWh3TVjuInEyni2k6CV2wa
hGzIO/PZutPd1ZPbDQoxa+XnCCHkRt7k8iOZJL21/ZbV44BVjhSjJ9vzI2nSOp41
rgmVrb1bfI0kNr+t6HiELLIKmlIDARHfyFaK0UwlDgh5Aeo8Wd2gcVUxucH38SgN
6f0u9ieq07RTjzWHCudIxYQwRl9wocSpoMI2bl5oAg5K/37MIgML5AQ+PQpBcLAX
Rvmem7jlPrcIoAqKr+Mm1EEzqXlIcc475Xk7pWD6tip5a3HKFciDRuaaONuAMNay
uD7mX5RRFicCOTG+FbgiNyGVbULFddh/fIa9WT4HCcMjDB6Lahsr4y8tHFNpZoXJ
lJnlyqfRjVgBiZ548gFOE+pL0+MtJwYQ6CZSlVlofEHM7AAjdE7bGwYHp1phVBJQ
hRDOwvg4yw8vKrJOu9TwxO4hC0NpAhA7N85WiIX4YnAwJ7xe1pn3b7Zl0h34aiKf
iUE1hRNhy0oUf9VCA2avcEu4YKIvUjUQ8JjIhE83exhR4YhDrmWnXwPzfS37jeeX
ObmQ60mYMEDLJqeYNhV4oIXFFSiX3WHdLOSFRCNDFh5paDzhXLhVeNZLl26tDHpR
Utto6ZDSdSpgn9TdJUijBadw7ZkBRC/MQvexV33gCuQpZXRYZtEKaBRLrPxA3BD6
CQ9gPZajLVY9P81vIOwmqbm0Opu6obrS85veWqmHzC3laCzEjHUEz30OSwUIbfD5
Te7+4r7Of29O9w3g4l3utP6g70f+MZ4cODDaRSc4rSikgp9qawpj/773NRi9/bJh
L9c3K6l/h19fgaVqIcj8Fym79snhH5toQvG2m/b2itil7Cs60NGSM55CV/pAG5Qw
X4R3srMnYKaNVniqq660NtT/TZ6MDzmcPm9FJSKsJDDAsdPHH4tW8VI7vvtpS/y6
ycRy7ulP0QpkuvPT9YWJ15JjE7FtZobM4IwnPoxyODRXIs1oNF/MIzMztdN1VPpi
Yv+ZY+adHCxi4i24KtDN+F4lL3NBe8JPKC+lbmXait/t5KzYbiTL03qTMBalQDGR
/APVfhIbt3B7CvswFZo/DS6dICYHBYQhtd+HEzQiNCtgVeQ2xVvug5dO1TwsWbEq
+bO2C/5h+GpK/gQHo2brdexNAO9kbPHhg+GtJTXWsUQwXuyJV0Y4dLTNgKIdvQSx
5qemBuP4sCghjRb1+AG+ygZzqmK4ySpym/n98zLxVrWkmCeA+oQInd4R26wORm9Y
G7fCh3HB0Do4tEV6295izTWL9AqAQ2DgUGkMYgS5GvwOU7mZ+vtPQaS4pXCSqwyW
LORGLH86IbCYyA4wcGznYG8c5cbv6OMcLEeC3I87eE+OdA/6+LdGQGTNfLI7j133
eknLvBd5axMcENxt+hnLGPGSaleljAVqrvQM5/ndywuJkbwLDuNSuGalXpnUuuBS
Hv/Ur8TngbtDpHaimdZjFmg8KgeOUqxgfovynYS6phDd5pbINoPLE5snPK77dyWm
2r8BtOxprR37v9uizKsoPQ0dXH+qoPx//ICefQTHfrBlermc6HsyF+SMlAmWhkzw
LrclK7Tgqlg8+ZIUxNQCusGPQ2rm8w7CMJ9j4ooVO4vTpcbWJOXhtP+XcnP+byOM
KWUzpCGw/0ECaGRHba12CffCgmr3p5aGcHKLa6jqVumzFvaFLiKogZ4p+R1qxgBX
JUKdUrR2zmGIpHnwCgrNzzdNicQGb5SI6JErxwDReOIpsoA97rwBp82ExoIQgoVG
9NjnXmceCiOjx9NoiduV5kWf40Ge5/iVEaVVjm0QRdjo/Ei+hBAQEgzEtU+mExrt
sd9q0xh8td8Li52pefRiRYlURCDhF4vHXVWoMelFANdv4tV+0oi4ELaqZrRefvC9
+zGNbcraehkJfev2Un14k+Q5pSV73YoGDF8zHUI9vVNmjKMV1OEFLhEvAAa5CxXK
yNCroCXrJzQAjfYL6+WU9YCkwC2AUt+3BzvtQ1jYLeW69M3NbR/qq7ir8rlLN+4M
a1h71QvD/qWCrHwB/8yNt3ouHXbXAIgi8nNd9PHTdSpw2V3Jvk4FXQec94RHb11G
URmBGdi5S4oaJRbCE/VWjfUTM+1jKOGDR0E7sWWUuuaqsMqSMLUgB1hxeGTWHAfl
8J6AaKp/gaHLt3V7dMhYW99jq4mkO7Nbi/4j7BMAwkRfsC7PFrkYL3mekkoepSQX
kR7lqu4ba6jCudFrYkm3KbTa4OUTRTu0RqrTJIwIV5eE7NCA9xXfR/6cy95n02Cb
Bv5O+0lu8RXSyN5rxrEJLpLjQAxGRKiwHvpdBcGeG1SVvicFpwQtMCWBTcaRa7lD
nUI+7n5BaslavPs8TFCswbM3HPiV1vL3MbFS1+x5Gew93wq8KGh11smIUQcf5ZSL
JdbXrJMHKIQzNbzfzj767gWeUhaHPTibF+yB9in1JhPG140kTZ4G7QyjxgjbL9Cx
TjXEJrAn/WmlLE2+GB78yXUc4QR21ZMBzlSiVgcWcr0MwsZMonIKYgFFFDyiLNS5
Bw/kxdKcTMRC42arAzSI6IFkuW4X9xNBKgy5JBf700jhkDuWKpNIUhTJX8HIUQLv
pk07WUzmG5dekrjuYh9CYe4UlfCL9xkZgIBVlOstOPl1lV9M5S8fvlrlJo2JrReS
O8t6qDMl/L2zvgiFJTdx47Ta6eMXMulVMDWApyrVDuvWpCfXkmHQ2BnnvvZYr06Z
LsQcwmeNj+5MtoTaESpWjfruX1aS5/ITCPKc5WOETqDR0zjUQ8LQSeC/G/2T33/g
pZ3cdVOPdCDiK0VE34F8MiN+kQsW84X8/cT14rPa7Y5yUpxj2te4H1YtvlhKg/Kk
0T/luQLEZPaYyYVdpjc2Es5SIvXCoJbvAei61k9RplrH7nX2MBUUVkxk6OpSCvjl
h9oUG2/L0mIMySqoVRP97NHzkLc3iRoafvlZneYVBx4wBnpG0hqAhYR1B1tlChoZ
SqyF+k69oA7mWSf1kZPcKqRTAhEVzOBfAtxcLsxCopeil+bSU6/UKivCLSNOkhFr
AavuLtFyU4jB9lQWYgQXMrG6HVzmV+0jX6ytNx1wV4Mi2JQR2S3HQkQhI3bzVuKW
Wbm1Zhrzv90k8BtdUjFDKgqydN8GFgRJ/lU40TTUSgDABlpelWk8I3GgXqnr8kMS
TxPKcrvqoUDlLCe6KIcuvDUa8wxY90Bd7J9YElvej9Im1si6IN8xY08DmJC//8vV
FNaNyEbUL9h5t8G5owrVN7vZavrlAOd1Rlv3WoAs/RSSpKQqiGw1ttECdNj7rkDl
2gLrnG9/CeSbUSG6Z9CalmGKIGkrllSeEXZZMr0jPIzfYe+/AXGIpVT8m4OT2QgG
XVU5QwBLZQfcSPqeAIlOops9ifCjYXZKYzgZ8iKjJ0M4m1CeIJYvhmhii1t9jaHS
sFkuvU78T9x9mT3NUNjnaK3ot8rJxjEB2kqx9Dtd8fUJ8YpqXoS9NytMKKC2NvyJ
B/S6XIdfI/tunvybBTx1bB85cQY9wq5OkjS2lbocgzj0c357szi6/Dfwm4LPwgBH
RtwBhGWokj76fXfBp5Z28x85BwSfl2IIrBS8KNmEtJHp/L0VyQHXPNTT/TwIn2yG
uWaK1g5evckL1GA1jZzvUz5zkR9K4FqW+xb+cIzmhk3h39OIZ4Ve7YXzwn4TLRDt
0ly5Wsiko+fN8C/NOlGhLXVeD+Dh/3WwnTfu8sLC2OabM3vylfLIlKcLK/Sy+nw3
/nt8X/3siA9wQHduAqbFoIK/atCc1sZJ5Qkuq6Ql1mRlJz4geso8IUOKMDRRyQVd
O/2ddKCW5BDG/YWDEwSU8u3whY11T0+k0t9rZuytF4BvOON9HWP0wjO3aXYZ3acd
alSMDjMI710B3Jyqu31ey0nyi//wJGwfSAN3C2675/lbeCNOI1y0tI+J35i4RGNz
Ldg8sdhCJW8kW+FGtHvuPPQvoA/3lc7niGbzPD0l6+Flk3RK1ygGykCB7RHung3k
q3ohRKwooGZmIOELflWosHBW+yW3qsI/kqpGvSn7U6aqj6fQg7l9yYZvqhiHyOQ0
jhVTmlO8qgkYw0GSq8X4B+t3m/NrUKE3EzKjGlUVipQHNuOKBvOCEu49hd5D76Mz
g65wIo1yV6LTlOn5ASfAANiO0KDa3ceOyXOiRdSziCUQy3FcPEgllAPcID4gqBpG
kbUGXEyfLmO4Wj8Zme51VvvtaNnLPHuXVm6o0OEtDdpySd0Hvo1TtSnesNaJHm0F
9dYZTk8H3XleJ8D2SlYcgpHY3C/kvh2DECi/7K1SNUdtEP6mR6QyJNYgujJd8z9L
OEZxWCjxBsqs0eQ11M2cYK7+lNbYRyRTNIdCciJzeWUUoRe8teR6b/vWiHxwf3U9
n+JktbEmyy95bp8Y8TTNC5And/j/jTaCZO4lhzdI+QTkJ8KkH7xSDAJvIGYPXZ+G
4yzDOxrRYTZKo8cSFEpxukYG2N2t9AjOmkCWgs+jOv0T6PWia23CzMO23JFdfJBn
GZ75kU3GXuNhDKyc9TGav244QjZHpfFeLMTvfCWFOARleoXFnNR6mBzwIrhJ43dj
kOzLPDSvpk9lKQgTo9CtYssvQv060OoNQYPkCcU522IrFShmDz79YNxjHQjibSF7
1QAbjeVRaNOlT2iWAwjY1c3V+qB16CpvoMfjjN7WyIHA4sNUYXrXdxYyQL8sT1i1
V9R5CCzjbQQGVBzT1OkHimnM7hcP9rLpQOGyH09Ic82fOl9tb4m/QWLU5Zh+uNZ+
bsS0nRfd//jBvMsjM3LcSu6RKFA1YlIV6MycIDb1ZbNDzZbNfHsv5k5vc789mBqB
6d5Jdgq0bB4cc3wC4IG3A2i/wBLHsQr6gweEfKv02be4RV+sqqOsDxddLAWVHMcY
Zwtv8lHJ5w+GiexhYnPEWoODYDh2P9tYf2i6ry66luh9Recauuxp3GsR/xzb94UK
L/RlobKbc5fULuv+4CO6M7VPTIaTNJ6HiSVjyctJPrIX13oFK0Ps7nQ8suJvvid+
Bf8hZnML0ILqdHlJmzXzPkpj6JVp2CoH+UnOyHQDcqHfUbR9RuBKOGTZ4xRtIhiX
Ki/nhZJyXHa2Vutw5Cwjiw8wqYgPH64w9zpC5lUX8jryD8RSpXxRKa4WvgtZrkMA
0SAWdiUTd1DT/0SpkxxthFZwoGwfbzvHKzNpIafFcyx/YnZB2PP9XvrpPQ7XApwZ
pnu5FQSHlbgCPdwAyAKnr4hPPDN4JPWmUAIOAIFV03oQtQBPXuYY9lDfgTOIdja4
dNiKW9BGdWKEbR6KQafL0jtxO2g/iQ+QzhdjsgfTg/Sqt6S8Lww+ZuqmcXzCJa/n
Mx+9IiKQQ4zY3J0ap0K14KU2xK88X6ZMEPxv34Uj7k/XMnsgdsgS5zQPuDccJxcd
Nn4gW3JbCsfpojTgfLIV/ZuCrQ+YqnHCqVIZI9NySQavomi0McNCGTni2yQkTMMb
6Xxl1J/TPRRbcfDfmbVpkw1dTun+fn2sZWunZkdwql2mXPHhaS0OsaRWULsDhvkl
PRXN+KEZJdv2yIZ72cZjdLFODH6xSW6TvJn5ZWjeV0SeGK/hIZd7lYiEDdK9EZBG
XAxUChiuXLAtZTtkkezVyp2cJgPo5PmJWjtpns/O8MuGknN5lHUlpaKznusZujYy
QRLuE+L6Ks4HFmQUh9wtR6n3Df7julg6p5iJvkk6OdDfRQn0zqLFgRRwhj/FyZI0
Axw25E+oWjkLCRFdGFoCE0BoLzegal9kY9qrHlDeLkgMpgQfUDAmb9xU+ZS/Xrcv
ytWkkAhJjVqiVlzv4/sL/0zfehWDOdmhY3bheqMrMeStZtTU+g2ILgD+dBfuLvF9
5jTqKDwQKEexy8/uLFHxSQxaLFqmBi6J6t+VBp056/W9O41w7BX2V+lACOCHsZQI
/A9I8b1AuqrksngTiuPtIz0NIctEBJYyCVyZF4bfCcaFAmtdvmz/wtiOSFtOGJB4
w2pfPbsoCDgsS6w1ZDyMdNV+H6bq4aypcNCG424czHB7veImHqfOclzqfItSpDWv
K3tw+gVRIk65BMVoqZgWUW9S51sqBxFDLBYWPQLrqJLgA+fH2pAzXD4yCq/xsZk0
NOiKkvqPvctAp3WZRfHGWxoM0wP7z+VtR90a2aIQTXTpntx6AUtFWAQD8KR6lT69
KHKQ1rJNAQq/euAGEaNANkFE8Akx+O3x+GzUECWb2f7TuGy9HLEAJ0LfWOFCERj7
kCU/o1/2r4/B2xARoGLjglMdorEvMGZZ1Rjd1QFI4Nl4E8yI1eV+i3CvOL+mEOx+
zuaPy2W4jzj6tqhrplW8Z51njiTAz916pbrcBzHNFKBuBP5kgv4rQTUrHmWcTO6L
8c8qdod0KELpbueZSuxMHn4OVV3si49EsUxb3vGwTBpgaVjfV1xbqkQ+bOVKNd1w
QRR2ffJc7u2r4PSe6Ds6/eahuv4enNGPa6vN+zF+8mAo1tuHNRIkhlwuVX+JeR+2
HFc2yxHOuD8jAyT/WitD6L6RxqxOJOTShhI9LGmuh+CCz0gPmuce558X48kL01Dn
CAJpQLSSq++rc2m/WaEMVS69TAYDoo3Axl3tcqLZ1fyf60P0bFDnQLpDTb1N6Pti
tkIyLJv8mj4TqZmVOv8jRdTeHErogo+b+bOrQJfeLiMK+P/NKzwM/XTHitqNd6We
uZif8bWWNpvomkxwLKJ8DS0L58Q1+3yg/elA+DJl465bqz9y5cJYX4KUh5lRUeHW
BiqAAbqhEM2Lvm+hndHwjiUb2ShCiQd4OgSaO7uUSMCrjT8NG7Zrt45wPP/kM/fJ
booAk232TnWO4DNmDihRR/F9OBH84V6d/y3U2O+RZ1j47ksxhW1Uofeqwv2L2cFw
sR6lZagw/qy3A6zMNN7km3TWTXFSwkbuxfxwjWUrvT6K52OLPFaULWHzl4CHALU2
+Heo8FOB+d1K36QWC8llMJ0gKtiGlNuaz23R8wIAZyBBQVJq2sBSIgOy4ICpxyrl
miCZir7FCZULdWAUaQg/MwBt/6IgES+rdHzbb3KW4LqdDiyoHoE6h6p8M0WjmhdZ
BaPLVpSrLrUmeI+OUL6cWbfNNaSi19zOj5Zox5TcWDSMa4R0QXXcxaAutIxnmSs/
GFwRJyLd5OMXdyFaRZNnsZU9WJW9TdevuhiFX6kn0MS6l4A4bmAajMuyNJ8mHlQX
Wxq240Ty9ZNf6tcvrqLJwtm8UZZuyAadvWVqrc1109+H9Cf9SydTvHnfGTbCjcd4
HYr8RwsqA/pMK+aFcFWS1HxCp+RBIjpEtOWg3zceK9gdLlppSWY3foFNlOH4p+Jc
G5s1rzv9LOHqfN2ziVODgIAshrn4tB2VTn/FS9bdR3nZ7xQhEszj9S2OZ/LF/Roc
tAK1gBMWr16YJumoXLzyYibYufPB/RCrvMFUkPcxS/36iGVwhRSOz0gp67KnX2VI
CRgq+U/GYbstEO8m12yydKLV5oZFs2e2sJxlnaJfqUuVRuexa0nlfh8iDv0QMqt1
6QEDFxfqmK/VohoGesIoPPkMB+0Vu/ufbYFga94yi53NHeAp9Nfpt4jWY/6XZWko
dAFuOIlLJTIq3nIjUvZMneYOOSMDJEasr040ESTSHdzCkUtj+j02skREVvJUW7+L
d/gysLNKJzX4NPOUllUY0xRCDHo0xYSdYKIXJcaYLerta4BQSrHI5ILr09bwtALb
v+QxT3Dz/D81dJ5goB6pFduA+LQd9wFt2dasufrGZOt7HkcfNaR+SwxD6tuMZ3O5
es9+2wzukgqMGvpSSlm3cgM3S7H8HVwJ/kgnG0T2OmmNs5I69odQKktTHWytBWAF
N/dGfuqVoAF49qQFvXwUGElPLb2wB62dwju6c7/Tr6CG0DzrMqbHpFRQtfMhvd37
HTW3sDaNUBKJEYFkKfiJnSb59EjAeVqhizIla6xk9Qh15slH7Fov8z4lpandVlzx
vWiJxTTmuo8XLKeXnkzpWodWzJ1hyAxizOKSfKvmCp4jqKOySRXbNWrdl8zUx5P2
CzQ4eVHiLrC7Tryb31FRqmQjnZRV1M4QXx0RNiA2jZ12y9+gD2oIPDFv5bD2dESr
lkz9+ZyfjP+KFOCR/7SR6IqE/1aResXrNvTU0ChJpSqbUuEQE1Jvdhgw+8OIIOC0
F8cE0SBcxG0VAx3iiJBrQJXCWwnudcXGGrBIQ3Z7L55mkWUsCt7bDVLGRwW7/CCF
M+Lg5ROyT8S1FuLOX3idJkq2WGjCmYSUIFEuYpFE+4wj7EW/ujuCL7kH7KpozukI
/TS1RurOrkdrtUQl5VWskRHV0B2NUjFZRzQdqIrIO+neeUzK9kMPoVxPkYsBTh75
lfGTaf3F1G73PLbBRyUTQwqgsoS1F3A2PEiCFEtG6tBrNB1UhtwBHIRT4CdZZ+Y1
HHvwcKWPlim2lj6vcTqUPFmR9ELFxMWH9NOgVkah4hEKeylc7sNw0zw2wuSBp6Qr
WcFtrLNvqDVAFd9dW1eN4vfTQ9FF5We0HggYNxZAfb/6SQpNwKCqmTigQlRwZ14U
Mzst1cYy16TFkjA/9Y8Admc6uKiLpStBf+T+7QohLzKXUq1bQITvUsQzouCjGVa9
HBAjuuOlh5PvbxzCETUd+1d9RLu6WGbwaybeb9N5K693VRbiVzSzJE/uDCNaIP4w
PGyoeTiN3P5aUp9u+VDkItnls6Hi96WFxKL7iGFIzjTwh5wElrSG9oMJDxVV/oRk
NwrfnzxSUxbIPfC1ROkTQrm+CQxhUIWHxYEW6sFpMcN2XmrGBacfA/EX+ByKUex1
tqn5qZ3Ru6YJrwSJJUm+SIX1PDzDlY0V4vtCh5AkovgD7tL+AptgpYzuWD8kaC0D
Idw+VKlSJx3RzRxq6uw2OlIK659aReH/M+3eKIWUgjeq1xTcxSyLZc+wrhOvu9rz
rc+V0TfXfgmQS3UcroBQk1mRchfzPaSrw6ckpuaZkh2PvhJiNd7xSNIU2GIAWXxE
mtdWKSAyyl9yHWgYoiKrgbqkFJaguE8vdWsfyO45uyQZQLVszHkwAnSxpnGrJMvw
J03tvWwcCXCwGUIPeJ/zHT+Y8lf7N7wf0gCXfbAv975Z7z8IUoGzpZhsy5zgw+A5
SkWVMnF2Tzi+r3DjbzosW7EIjGYkQne/b4guio+qDxTWCR4Klst3CEvjOeKuEpIp
fL/RnGsyUu1UyBCTeztjk60yU8GAzcZWaiSDJZwGbbReRc9dY5S3aZ8h1JGCR+V7
YyDorqm4TNl+r2Ho61ORxgN5TUfdXknb2v6UIN1HuwdSiU6kAjMUL+ffnUJ2tu8R
UnhwShfEz4kq4rJfd0k+rR1yt0TyIQfbYemtrji0zkKk/Hp75yahUBpzqnJFxMmK
LMmwAnpv5q5+8bDNbMETOD6aTmdI4R5QKtcqz9X0h/R+8rAs2Hm+JlRRGuWSkEKM
KrAUY9cJ4my4Ehx8Pr8unQlTFYOiz6FYb4ivTPTDtlCqoWjkHDugphLxJ24ohghV
NQtohIayDx2NNAQ2vRE299eXb+nJMdq9SSMT1SaBLEdDtHAW9QZlwaxEswW+MzSF
KLPlk/9CizVvFYhdukdfdy2G9RD+T10CqFtFbgVzHqAJdzDk/BwLe6ns5NLUMDf3
ezLnW88ndrcs7EsnxUzJYqkQ02bW2jtsWfjcZ56yax7/6BngVOCCk1ndU7Zz5Gxo
RICeHSWmCwEcBxxCbDbQnbI+8NF6gedwm/Bis5uFL4X5bokPZdPzO1G2mUOJDVLY
GA4x604c5INU8nEvA6oZ+WNmIQ37znKLtMOj0fVwB/3uIPnUNfRUPxJUazDxBWtz
BeVQa2XZq2jGvwXp2Q8oa0qhrVH8Vx3fz/9MGckdbamVOQFc7++9MGTdgE99tv9z
GkOACPyBA6EoPBbhLeo+/nxtsstwGKyzGuZozP1Xqu5+eSwBFqOPBZ9ckgt7bA6N
nT1v1NgV7I3Z/Zp5jXtYqk348SUJulUHVipmbX/itSu15oUjvaeWp87vqXVu/JW8
3582I37dwUKpPcru8bv07toOjfliHUjpirzn6Yx3JGP7VMJDsIACnhOMAOIKZnxW
sBUrcJ/PDU5wi0/5d25yiR7OqU7xu8ajLEVrR6CKLqkPeeYFWnIl0nk3qraj3RjQ
cuEsdmeNxGTX2sS336dqDBgqELbwjdYptEmLiTXhEERyJZI61yF5Ub2xkfKuRdWj
IAht/eso4HIhJhPoHp/bYGRi6h26jR9UUD1ok/Wcl4ZYWXv9obkmMnRxhPBzygY+
YBH8XiLaEV0+weINVoeuhFslw/9DwVpcvgKHH5VaB1j+j+ATGuoy3jhTODCMO35t
HTpKauE/S/6e1lxkn4yjXNyRm8p5qioSfdTOfABmVNB4q23r5VpiuliSMg8LF8b0
dUCM3iL3e/l27GEHx6VsuaKgAIWrCTyGgMIyUiEGdYmFKMEIXyegQw9YD993gse0
QLT0ErY5xx67BFjL4BPdooGFnptfUGP//L6tFAi1NoOlfjwlu8BcCnSsweHGNPDr
JGwyoy7OhZX4BKZzFKrEzxXoQon9bIFHv7OUwIyUfV9yzru/nRttbfgjeTlvsLRM
TmsvJM0MkpIDKOK5Szr8LpxDX5Urcr+JlrbD1PAWuwOLud5M4CjHoty2A2hNJDh7
eLcVjMoX8EPFs5SyQfUDLxiPPumlSGeCU5rPJoy3ajQW4NBKt61DN5kML5iWIEA3
O8cVvNafuY1TB50Wt4uDVXT6iQdDxpgfeq+wWrrbmk4zkumfgd7iTS+Q+Vft2mat
zS5VXnvgI+jUMKejVwsdHwrX13h85T70QJUV2aEp3HytOt3GT4dvODW1zLaX0Hvu
xAUKkGzVGdqX2u04cjKB81IzX1u5u17iDvYRDQFi0ZMViS+qk7LHlN1Yy8/+7Mex
dG3w/Uf75YXuUyUVJ5zZtjMR1gE9vtIDNmQ+2P5NLS0Yg5Wvb2ta9sinDbInVrr2
77h/699j9JZx83nEU0SuhTBkvCVkMND5Wq5/dCVopLzqSiHZPDvPQV1RB3WnWCPi
F7zjdY9TUyFLfpcaomJjSk1qYfHUhzh/O9UIdlLQoXPH+H2XhZdGJ/XZ10rV3GE1
rTpcZA/B4Mc1u9NMNJV2k9VzJlhOtwtBEWYlKF3dYuwzjy3ATc7xsChzIxEEX5qY
shKE4Roi4TUuNBaqoIOEHg2MiDVqOkcUDvVfZq/r4bSBikCe4fRzGIAS708EVXmH
+P3kAk+c/hRyMyeNa674eSbjnwGBmQ76wd/KLzww9Ah8CYkpQaXmlY4MFopV2gIe
PM8iAUbZI2yxmB73GEMYwa1mcOLGikiO3S3gbz/HOTP6P/RqMLk4x6z3qY2pq9Kn
n86pRX8mkbEWwertpMDJBhU9hVkj1GhVRo5Q4oeZqpyO7Bhvhq/WJd010luVnsxI
/w4xMHlW/tqCRJq7xXdFKuUC1tT5f3L1FyZSvOFAysfQseqEd2it7ljKIasptI4f
9uUAYlvwaO9FcIT8CKj+E1DBc3sCooauGiC+hyPzoFtcrtwio7DjRtA7nWYUOfAg
IWjTo3Zvn9vDlk/pMBA5L7FlciulRNRCK/cSIoRM8cNHHPmWCz8ERN+uvgf8yJJ/
oLkjziWMz/hwJpEohalgHG+s2UL08lvM9ryy2HnoJQQ3FMbusiWRdWXolOznqeFI
uj2h6uQ3utO7334LaGFhANm8NpublnW3uvozW3WaXHbvuMH/wX7tBsTWB7daRWuV
wUzxrrjOCklGNcgBWrih8rikGJlCheZ2empSebeJg1LcUmmgY5IdGyg1cNoJIolV
kEe1miUdYeeBElO0RjRJB0rTYEOZh/Aj/3lmpPM6rolt4x3ohk7dyrP88YIVOAG4
e7sYomisiU0tZcVtDVgrLwgR1MoJF9nbrVGrcDw4C8F1IIy5bNro2aaRUDW5p6JR
cA1S3J7Hyp/ZqZfz5N+imG/IYNcn9Sp1qhDCwzlpOsMS0Hxn348l0KVqqz6Q+X7B
zLWpdrekJ9SkXw0G8LMilEYnYegDoLSMEp09uJkdfw7m1FQe38GOahmctdB3y3gO
UI8l1f6aD8LpqMlBu9vB2pZi97c3WWOo8cWvszqoUqW1BYpgIjYFHLdhex8BDr2Q
XGzeLWITvkhpDOaIMwElpGGeRe/iId0ImBiEyDX8/aKRALa/kDscjHYN51M13n6z
wHQK6oL8w9HV5K7nmp/ZsTBZERHIb2zlzteVyBU7XH7sI5B8GbBvjQnK95U+hnML
Ejk4vcj9uMwj6w8qlYz2l79fk7/fIVxyUMWi9kJXBzxnAJNxBAimVZwrCJXpRMF0
/d84EHShAisX1ZtfGlgTVLB5otQ7Z/Rky0Dn2XvIEBupybGItREz0O5LlMP+kI2E
p66BoU5KbWRFNozVP90NbR7u2Hk8cHCkDWSN6pH6vFdUv8dWwlnBnHfQEPM3QGIa
9pB+RxfIdsmxVQxw+99FiNQYNnkqoqLEwBOXfHQu4rU6TgxU+g5oVP3tJg2tVUAd
xDiiF1fcajV+ze7KYMkIHbFfjtTTXP5gyMAFSLaRtNDbfpS3CVDPHMiNLIdcf+CD
Z146Vb1jIrb2oDWPuiebkn5nzLPvnw3K+zTWGwfFS+II+bhDl0E2noFoM7vTiM/x
4ooGYOsLLvpjoAbizbAxzfISjrTyZeTVo7j7+UJX9sQPF9TKp6o0fVSKINN5dy9H
Gk7pYQPw11fhqlP+w+LQSVpjXGTEUuoASDve5O/02nbWf9HbkCnMamkIxVtwYzcp
LPuBRVag2bUu2n/DgXO1TjvMW01KqCMhqtGsHAR7901FF9yc6josu668PlXpEx+Z
SrVus3wS1Yp0KwaVjfLg01lE11hNNCkh9yjO/gQvgEjaY7TXV2sHB2LvsgdIrrBK
FV1UsGM1t+RPx+HQ1ZtWjEkRyB/ZW0VgM80dpSp0rozDfsMnCK1uysddh5jw8BTB
mK0RhdVBsFhSRjEnSBDycfODY279zy7xeIY7aQKyiO1l6g02E81+7noCTnHIy+vv
2ry2+BJotOZCV3m4swfq+Om7I0wKhQaN0oggic4feM5S0nhvg1HlOYXjjy3tvl4I
cOHiJGAAiYFGLwFEbxD1TgrNxdQayWXWv3OGBJPwRTSgdsrQI0pQMpKqeOQJn0T8
++Im/CJ5wABLHre8LBcUNzaCEfhu4mcQQBelajHTwdeD+wbcoPHcrvUnq1R/un79
vE3q9WhSwUNyT1jtA5aP5BmTBa2NOwMgOxSV7RkS7yMPWt6oStrkk8eh4A5AUanm
jwTXJMaigCIaUXXsaVj3aP22jSlBJL1QiIsyJOjK21vfcB+e9G95i5fW+Xdw4+N4
343uCrS4p0Nq3JY3qMtljByiKTCmtrTpvB/eYukYqoltBmuoG1pLqVlGlgEklEYT
9ms/9qqhuN8JaAJlpotLMNf18LgkHCUyoZ78MBySkXhRs/sPFsWVx0Y0qyftGk9Y
nT5r4LL3xKZBb5im44yuecfI/Z/ltiWfUt2dXbQdq4NaledPOSgeQkDKATS5mxtn
T2lZY3nisWbdp6H7uqTPSx/PIuATUQqIWzfJGGq83eBzuVnbI8ViQgbaq20xkyQE
R6TyegNuTYkGDxNLg7H/upf3ME4yM+TnOPMxxEEhyfK7BrTstxqYLrIO5uGaHNlC
GSzt8EKid3YYmCoszuJKLZOhilbXzbgZgWLy73ZwexH+VCopfriJPcUaKFKSL9IZ
tN54B7ozw0dFT/ksCsT3RE3iljxRIYs/ilVJeRcWpr68eOFesYvGrFoMmbaOhtyd
dIhr8ghdcheU/k2YUQfWZkjHDpvcyzbIRKoCG+o7aQ5RK2P53u2Iopk8MXNeYClf
dQmZzdlPmIXQjdexSHXXQSj9Ek0jDPhnVml+jyw6ZWAvyIkqn7s0EqB3nUHliFSO
M8dTcbxB0D6MLX7KPStCFO7f2pm3DEZcNInQ92fgGLKkLdU/JBTKh4Bzr5tLCWTC
ghDMaa8FvIUXY37hNaiKDL1+TMOInIHQAJCe2ustPn17d0fnRGLnG+nVceYKWdOV
Q8gtmQ1iFRQsdxzM0VA2rnsMB1Mcz8uG+i1v+NDryfxTcUyymrf4kpd4uOdpR4pR
VpM23aHmSjAv0VsPjoQN3fmEevtEvg7mh86e0Xh3CQ2w0ML94GUtTBc4F0kvEnBb
e1GkeskP3zECXsvx20fK/tO5ImlTjs/oY/PKpDl65SBL33/fVJZwYyx377oeBJWn
0mQ93702pbYBu4ao1jm/bxxXTARlL/OarKPZcLinQy0Z19Ibj50uAzh1RGvgyVzq
LIS8P2WsFQKvjBBCmGjXz1Kv25bxEosYSVPPETze2SvPRCL91MqJ2BAAdEMhbMlZ
gF7n1HR64Ruz+UiVM3wkihYTCoKk6/Te3g7zBnACT/TaSLb9TaVf+j0V9A2vGL1d
lDQepOfPABY/oseXyK8Jz37M05PiqfdMDIy/w9dXZcosrRULB/2tBt5lEwczo7PT
Lw9nE8hhuc553zsClXBQFTeoPlBmt2kJNtPTF0ukdu8lLPl/H8nCxjfcY8MUwgap
kscYeaOk03OF3BI0d6cH9+Q0JP/r4tIeSljrob5Ne2foIn3u6Zv5agCEly2Ouhtg
NWEWk9gx5fsmwXzHPTBaHHAAaxj8N0YZtc/ZX0IHScxGt926JfKoU5KMgu5NQvPq
xdsCIVBkkWZFG3wGsiUMY9ar8YX7PFnHsVGk2s56y4Y7bnSF+yhmPfdigE4TrGOT
H6R+pRtnuLb2VHv8829hnDBeRbDfa6xnVS4XBWIc9e8jzhhSJQ/Qwn6LyA2b3tZs
HxURqRHEFvlQTnZil4Pi0s2nuvQW3E+zpEIm/WIJcGwh+UcwXb2sGbdT5S44OS1B
Pn0YLEAtA+0Wtukv68JGbEWpQ7fxhk11EmcS2jTnhA4hZ595oFuvGKVILy4FQdwY
WexKRNxTsY1QC2AI+zSELrhXgYksJxTLpcuBHL2qYsOAqD/PvaF7LlWhsJF1jjC8
gDvSIAO5v5z6b3TahgNh5iLg7XVcX6SE9LKUW/MPu7us+qzMQL+pNGjW751NEtuE
LAcCAVGygDMcKiWrZdBycQATkR/fbwyVEaBby+5MJ4tbfp/e/PlN7aUKof6eEArK
ERB2ZBsk09YL2awN4uvltP80MszdvVOKhi81kv8wfGpU2aVcPeFa06/uUT33n9OO
WZiQH/bhW5quI5zEnJVCJdg+B0NOvothIcl1jNODgx0HhAuwJ4HP4dhE353C9S6B
aAgptRGQvo4mFMDVsp9opWc8aaBDjekEuBOiL2EA08O2WBZE7FAV3QLo6VYBn+4J
HItR1GWYjkFcWeZjWy8/UzZW1Uc6xRstJpqWKi36EC82sKajbZvDfpiXxGpCWJfD
R5/H9vjlUQ6BsodrhEsbSGbKjn/10k/gkY0/OcubDO8svVFRJF4/eqrKHWMqdn6J
gOvn5UnCxiEL9keMQMQShiDj2Fwuk7VcS69CeD+W/diKo/TMUeifrzWLRocaNYRk
Wqrcegjq8dVouYzIUX5pH8g8b1Zjq4VTVHAaDJEVsc4nf5ck4LtL/UEpZSm8glIR
ZsnVfNEtT527pg+8JEmLKeMDaQVHcXlL++2Q9k0/kbBODyj/FcP6FXwNwj2WjuHq
qEO4n1uTuPO4YquSywSgMfkGLgx5q9CxShybueL8FrmNYfuG/gAIiwDLsVHhm0lA
vkWMTXV6okfrZZBuWPdalv71I6vsyzXFcWSlkTwUgFdrnI5356x84pA/8TyYIhR0
TAga1aacDE7wd0sFAIbXn8HMcXznTHv4IaCeX03FLe7Hh12pa2rLaGIZXbAnoYxw
/A9/20ZA64FeyLqcOlwx10ZtMbcbF4tkaIAW0z3R1qXIC7gXWnXRzw5NOKoRV0LA
TjyLDwBoAaxmzvgRO+sXB3e6ijKgwblSOPZsRJDW+7R+jDaDmeaunByKfumBUEJw
BAz8KchM7/KHSsQUiTICvN3vzVpq67z4S63vt9+NbXlu6b5UaWPNbU6Wse2OEqnN
4liEXDU3stO2k9BJoeqNntEvADYn9Cn1r0/fwefJ1o1PJld9pEFrG5y4ZjbZX9rv
LA4ZkLnof33zNQ87X5tGlLwTbf/Ew8I3EWlr+JrKmV3ERbTW0Ab+lyxURDgQoAa8
huIdAQvFO/W3y8AQZ9H7/wys0XwOYMvr8ygjE86MYdQ1fCsHIL1hfqDzkRMwcIFR
o/4QfBckcFaUnvdeGCs3Ih1eCqIHCaYBFDMh0DZQOdW/z6W+lJneE+6gQho4PWsW
1rWWzb23cq3frPEl1nl9WQrkhLmc+BroE08bvTVr7riY4sv/ROHTzJX85coAqK5I
UFdpLa6nRJo0nWEeu6qKA0NkFct71lpcrVNajKyN+o5G5ZRiNYHeXxyjodD4mgW2
ZvEA5EssXJhoGEVAbBMSQDHt+24rTvPdD6jWI6sg3kQSaUeokn7JyWclTGx8hOyv
eNjlSQDS+YnAZoEPYQk+TZJZ2zt8ULAILFDVTuCg5s4LmzW+sjjt3c5PfxOl/9J/
x+msZjMzTzWuZhCeNH30Te22INVuqNrAh8kF8hTCOuLdriEF0Ak7CEbxHWzsQTtE
pszX3BYljSjKo5BTcVqCWeA0HkrHvmHHu51DXvOca7+lYj+Y2itDIU3OJRl/I1FP
zkPDwem0OdNMVJTjMH0bwBOILSDd4s/oNcGIcm/G1jpMvVDyYcWaK5fGNLk5DYy3
3vLcqWaMXk6HMkkW0iImA61jtvb8DDW9xmg1zlCfEvwjOeVG55Dtow5e6kau6QCo
HwZn9oStsXoPCH6EzMk/vcKe1uFztzTswipbMR2RME/WMBV2Na72kmACFWjZvPze
r0+W5x3mu8OdSnPJ6gk9W+eZGIYhwXfD3kmippPAsMASTOmpYW6J7tB/x+D0h1KK
vVu72/sO0kzvz/fhWFtQr3faEe600/3AgMF+P9beztoW6kOZuLr2uvBR+yrKk2ql
CzRhLHvP8/khACyCSeDNN8nkWulvxEkfaZESt+LAuGDvBF4iayruK25a6h/cXClD
Pz2q2HFQI9rDrFmWbHRcD2yS0oNPByXpMbXz7gkmO9Iom/4zKNoe+KLepmYWhstk
0qCiP6iDkwZ/RB6G2YmVIo1OXmNgtXlMzHEobzlFWl6XBc/sEshF+HNUJG+e+CqE
67glQVuVi1Vp+BuEHGZ/RS+8GZg0G3rq0AYAtguzPe0k/felnsVk7JykzmqWnifB
ihn86AVvIjfLL/G/5B8cODv3+piM9hd5b6JXLwEjcN49FNWB0TXnJ2kudZyC8jlz
1oekJvPrnCWxQtnIZHYbtlQS0ILf1mKvW279NBVfa3Qc7crhfBmhwQRos+tait43
YW72eAVVjxXm1PnBu83WfGLF3fJDl395adcf6g0vpJLzKjgYshXyPhRVCz2r7aq9
qRgGQYSb7R0wiHWtdaZXBQ3SjQAUk8MEtokqnaTElmuSZqXxYToRAuKsdzTDSnrl
TX+WBWgSg0MMvkxdbT2gmjVA72/8mJT6USf8zXIhVJr5srFBb4IhKp9DvXoM504g
ekhdQ8cCwD3b82DZ26P4pNZHKMiBq/nx/Ox8yPVDL5841GQI2v8X6dII5tOzdeRJ
mrTO5HCFNpXhE+KvmZo2j18WETUM67lTBnHjpkUD59WiFVKKuwXXEK0sRf7jVX+R
Dw5oJnM3or/XC7Z4q+tL7+vCjgL421Gsw6Buja9qzRG0CfYVH5WjK9ELVIMh3Ndl
BICwx8d4c69TjQLIpNww5ax9hVjTruup1ev+sVk1KJHHv1OUJM8+ijyG6C6a/SQU
v5idBu6hYgn48mv7HEDu1dGupVnvKJ7NcxOEEO6RICr+LYx90Um9wj8AftqIuHE3
W+mEldN9sQSELiTA0dfYdfwasRNThfVDyzLYfqZVlXKpEBMFmhcz9xhvbdCsXpsP
sKztXHP5fRmAA9x+0LLyFWIp/OLzfEJYetgbpPF+ee2cem5Efr0gyYistrWKhrHY
yps0vgb6ORk2Cz9V2zS4VPXr4GP4dC5he3lwRavZLYEgEPSfPejHZCR6bolCyDZU
Vt83yYf4CAHHwxEm74SO0pskY3chDYNPvYa7fzDS0SycHp3YF1Il2wUbxHhWVcO7
MZTriC3Lvs9ZyRdvPv7aXBhns4PgmGrxeRq2Bu78EE7fdE0Y3yyEiJd4gInWZr/b
OrgP1LAyPibEnUccAoUwN84JT2wWuq43hkYRJy74Nk83CrWwzFVwd0qhTDgOJo2L
yJle550XHFJ9Nre3Hk0oGF59F6jFGwMxPpJASq/LsrXiMvYUCIGEbE2KcgeJZwdP
J79otZhK4g6CyXjkUwv9vD0z7OpCaisL4iD+Gjzl4YYSD5Y/frX/BBSU3c9o4yhg
cN1vwWCFzpCON55bkVzAWlTIN8l1X+WcDL50oLAuadsDvDQbRzRiczU1ayY9f9eI
1NHtGlm0bnF/k3DPUd/QSUV8rR2jAoBpzVLxwHp7pedYBtty86tXyOEUGR0woufE
Nqxr9/qnslZ4XJ7Xry+WNW3KphvZOgJhPwiBDvKaP4mHnSrI0f2KJX/hov7MiHyw
+TCPHkJt41v0tY2mjrFJ6rpQZjdDkGd7bUKcPESvJmzGlDNHDQvu73fuo0YMqoWR
p/+XgQn2bSVnbFkqkJE6mP3IEU3EcIJCoOVV726+9qpxXoOoD4vlDbI6ePZhiIzo
9Ctls+JvVqZy5tgNUE2GoRiL9nOstuYkl9lqFGoZ++Y6/8hy1xZruDXwcIuprtvS
VcUlg0IxliSCbwiNah2g57qcWW/ot0vroWk0rYdE4fYaWPviutOTkcfRWjlM1QXj
a3uhxFfqKqLXIx1nflTrB6vMoy1LvPXYWsK4Kdw9F3f4sD7w6c8uw02YhmM4tgFj
FahDhuFW9Zmrk4Ryc+0uG5/qC4mNDR4uSWp1L8zs+WTC9nJVFIAiW1z9MmAhOq3p
SjKelCbWoccExPoSURVvuFbPN4L3ZE4x1q1dZhqEe3lwvqKLfoHKnPp1JGD5qI3z
5oP2WLS65mbqof0zfrHSsqUpxKJsaPD8kJjhWmGnElWU+rF9zEbX4Ucwu4gUWsil
4gsG5moAJSmYhDM876+jXXorKmEHOtV6vTs1W2JezMUcuDFRZnZzpUz6LzD11RSq
cv1Ghb2IpzaOG8q2UgFL5zDjQfZNrHCDnTZHCxKpQFNJpr1/qHE1hApVbg8vKE7x
KjEVxgzbrJYNIJMgXMTdn1W2EUzkTX+NYKbA7aPsenLzFIcPZRFb3uJ7Dn0eYh1Y
I41KJ7iBhcCB7n0nT9HgThk+F4KYPS1bgUJHDvUGmTKEUW9KcAx+VJgxr2zuKbjF
zi4ChG4y/ru5fKqIX5UsJaRTF3A9r7ifypG5qtge7pvlIlbbrth7ttYbdYHz4lFc
mrOe/psYloYrZd2cTugORYa33KH+kAsG6fNyWFvPILhbuiLVqMdhuU/62gZPnHkR
Qwbq0il0ESLfdxEu4X1+REoHfdDnPSLYppnuxgRRGjqN+JLOr6XMZKCCuV2Qnu3j
ptXrSBAlQS/9kY3hKJsq3HNobCoVT5jaKldM7t0Ebs2NVKobUbEWZUQCJFWUH9+N
CNdW9ur+cIoaVNxglEh4071udYOm1UtvAvFK6K5HwCae/0p2cw87xLuptXIZ7D6u
UksurwxvqfCCrvEXIb+M+6Vk0xnsJFFMMZqmzntBm5nJOez/m6pz3F9275Y/2k2y
YQCXlh7Zowdcl6dElbGtwWjYunsEmxyUrCyVpWzcMWRlE+2Lrpm6P+B0rOZMUfBK
2WEYidgZzNb5IYrUd9C8Lr7DSSfRKPP/Dq6L4izg93Onb2RBUxPDL7L8pToxHQ/K
ptc3QG8t/kEcDT0xUwsgvR1obBiDaL/XjB7WJqdf3bbYymO0Kll65HqqqENWxoYU
ZxwYune0O+hS9TC3ZtY+WLbH6S3bjFTqMkPQ7Kv/YGTyQtPeU7zQwU3lLjXzfN9v
Xc2GLxfz2nFFUCgkSkfMb4MlMOsIYhQiVPE4ZfYYizgENMF8I5GHxNlVAJZX6Dku
1uIr8rK87MWW9YC/qWuffDiYMmANBYFmmBD/lcQyFUg5i+zKEVReHH9ntRRDW1iK
Zm9BUX9BFlvBS/mVCXvhTPN1PEGID+tusPjgLMptFKjGyO9sPfZ/3XJNAaDxRftD
UCABJkQvtSnIEPiTlQklLpiZohy5keY2w5AKg6Sc5j0jpae3V6IGaF1C2eNtLOSA
sCV8YAsqKqNeHWOBkGYdVoFB716ZGH3/Kg0w5RPbzzyXsSh40bVTvVzTwbUc/M4r
rZ1XTU/mIkhaObfQEqdl6s5nZaIXKFcji3BaBrzgqCeHO83HNozmltiILf01bpus
xDfr+HWxFRyLl7569bcY0nHgcxIRK9QDrSgLVsD/TEm4S7xCvVi+6zAXINSkZfNV
vTxjxB4J6MmdJOVWQCArgAH0ys7DObvff4/y0+8HhSmGb3kZBSCTXDWhP42Z1S3T
hG4Mn4UKKLqL67/1LBO/jX4GGugRbA0WK0l98bZ45ULQSgbWrlJoYl1Y1cuKJBd+
h9cz13nhy15WRDCFBek9nt80io4E3G3X9xpKaY9tldhJB4i8lat2ycCoOyLawbGh
pQD6U7SZ/O2689HNboAhpDf4shl9wNskcPll2CSwafXM97ZLjadcFPTwl0dfC6LV
oVdvApXXIC/EUPBBWGBsNVoGlldTYyAefmc0OYKvMbzVhuF34LeePgMqGuR2fybZ
F8KyTjuIiKTx4/65zaTgfNh/UCwmapNGdlkqCFL4lUyi3WzFKpqZC2WxdYT7+GaZ
P3mEhwBRTAskog+/Z0x4P1WVfoWr/UJB3bECkrCQ4hf89fXijHN4FItvr7ouTY86
aGKZS3LSYM6FjPHkvBUp5Gwa1wxwevCZUR6AiScSnw2v3/e5vIH6cUW9zLlTYavz
asClTLe613Ywa0epuT7tBbn5syVw4Sg73HPoWJCXtDFhr7jk8xQ6Bivc7JfB/J18
vinpQSh5a9+i8uwSz13PuqjbASz4gJaWrdLBdfeaFvHG8K2Xqo2u8LNQPpKASbkb
oe1J3J4kAjFLleL590u5rZwLfrMG9yHk40dErMbNMaXEFD0K2IeR+DiQyKUlKyx6
fLv7CcFp+kgYa+o4XrZhnjjOZIfhzWxpW3YE0oepSc/QYHIlyzsQiG8BmRkGBcdH
/zbyXq41WLJaih4gZPFEVg2vj3tNSnJG0tUI1gUzWB18kruXbVtXVIJGXn92GLeu
rRHl3ECOpJ0nmm1p8ZJ7vgSMKLl3Zno/9cX+h9QIVSts0bwjP6MY7LvrzFBYYxVr
2hJW5OiahX75RJWiQE9uqQB19EMQ61Cy7POBL/n6XMsyxTYMv07u+CY/RfNk43Bs
lnOEBXCnDyAnL3dKs4MIgO+7jAR/jHgbPsmrZPk3/SbkfRhfGoXg81hhLKPHGKAc
+qTH3sU0Fh6nCMdAXJs8MKF6vJvIrl+4AkQ2SAYsbKgQOggczbE9uJ7UUoVAt7FW
QkiR4ruSpmxRTfdiq8u2W2oEu3G2fUCtDtZ3DqZcjBss+JamcXyBKrXWl1LckI15
sPmd1vTWyXZ4yG+0X9RYn0atGuROIqdRswGbvsR3k3j2EgPQ+NW9ulY0yaeoZUNQ
NhhdA81hMeBCjrh63buTgtcyP5Z+CLXyOUPAbaBFUcZcdj4eOsialuGcB9V6Cdqq
t5TAytG2xcropzCHMVE4cenwdA7XcgBTI5pF/i3bsuuj2N5fzcGKIoEiS0x4ooXu
fJP1s6QQ9yYuWFpLOotgknd8Lz2SOLe2ie9y3xjdjavjf19q07gSPQ48Tp9hWcm/
rnazZ/DBhhxvICeSdii401++x5FloyDuQS0VxRWOcuIx/zP9gI7cgdIBCUvyUaJP
YDCWf71C1H6jP7R2xvnVRZ93T6urDeb2q0Xyl37o1F1+04nsavoK7tvv6h0k+XFj
br1UGClS72JlxZjeRdmoqNz4EW9/8HWHKevTydXwFlI8Io40Ug5XihWPEPBqzose
kPzqjsEwhNLXOTN/cjdnvDUbNQuwFtG9kCGsiv7q56WCJm9O8V7HFuytqMlSluep
xy6O4Kg5eFNfzfNmi2RRVbM9HqWvr55xhAt26sAfLzHKILWz4dbSiUxPZDTodze6
QjO9r3jvd6iEKZ9vUfJup08YLMUsMPDI1jLSTorhIWXwVqzfvlhO6V74qZaqHGmX
SD5k6jJC3shLMvHvGmZyuFLMRcPJ5vXA5QjXUVJ2yRIPfBf8mV3tpyb5wlcF9udP
wgxMZytVokvnWiH6Brms5WrtLueiSkFkumhIRYRCoCshaf8M94YO5wcq59kcN/6I
pskSoX74YfWCJBMPRRpSisktPzHrJpQWjL97oVSbsDMbmwkbgRinPLONoE/UZ2Y1
F6LAeojtuotYXbeOS/gAynuGTflVVDUDIZvVzqVykJ0YX2guvkAk1kvM8d62vg91
8sio8ZlqOjhjoXKfnhGSECpS8TMYBaIix7ubWLlWLxuaXXRwG3ze1Z4CzEVRfyoo
xTiTdQwJjO61x0IUaOLbEIlpZ1tHCItsRPQx2hPNupVR2YaujJPQIsZcMLKK5ve+
pVbZxv72+Wkm+DqnapEAcsgOII99Uf2JARiP7j7g1kNM8XAV4ebEOib26NY0GQ8f
yltX8eN2fp2wvDf/gW0Miecdr68pkZOBJ4dx87aekQ3NtKqUH3XRW465s0a9mMts
NwPLwUiBKHPfbt6aZtTzYsJlibMOjZ6Vs1ViA6TpQevRssr+nqXHMCeEICRqDd4H
aBU+ubOueXMPPKtdQO8B4rI+OsC1Nh08c5X6kykDiBjrx6W3YN+46UoHFgmxiRCL
rdQxS5UPdNxpAdA1Th3izNvsgA43YKymomtVEmsf6YPxpGCVO1LWwb9XOgyjF6CZ
1tnF9mlQrBkeAkB3Ax14COS/4jDibMoSuy9F1WA0octv+BKCxWpXorM03lR8mRoe
kQCtd1Mk2jQbBjC/lNKaok5hE5sIjTRihPN8vrMbwpYp6cvBHg4KjQxtpS163Stw
ZUz4J6w9mqplCNbr0bun4FxP48pmGPQE6wHzPjSVJ8fWs2SfTRULD3zBuH7Sjg3q
MNvMZhVQXhcUhFaSKuZohJ56jL/YRUoR4TJbUOEE8lnVBX34sZIh5CTnjPi1JqSs
5b8JzzeMD6z/nBAZXvtqOFpx/2jzdND8e4TjZ9SlfphLoJ3wPZv2XaKuCIt1XqZm
qLNFSyaJq392b/s+aHhC/vBD3PWu+N7VilCGcCK1SNzNMAPhDLGRHmWDpyQkU1n6
e6LqB7ND0xMgwpfUm/SIRr+MsFR4nAYql0v6r6maCM90yT7gMtV1i5rtO1NYzPSM
wgmYihOWdQheCQvBzPq2X73IRBygohJbla0cHRns2gCu5d0chS9vkG+y1PjK971f
BQPkDjNg1/5bGsC7LaB/jindazvPWmU8ctVUQvz8e5WnNATxBRtpWuvzJ9oyueHc
6IbQuxqfeVxaju56jZufQMdMmtwiJNKLxiGskC34OdRRL0VPNvhwzZZddXRRSvug
SuO7RfNgBekUcoLY5SLtaYBKQNN0/xzdzXI4L4RFV6adRPbFn0Xvgi7KJHR9toU3
zNOYeklmfCLdXb2jUTTjl7Dt7U86cBjgEBj1CX3SP5tNTQA3B7lusi1FSp+lQt4v
AQp/ecYENv3B9qS2avqGg70/DuJGMDsEFCS7CgtRnTrpYwkjF6fLkNzrnnXCu4Ur
2wSYSrACKOLF7q/0iI4zfxKwfhXDbBHdGJLXXgW/5s1pMvFHfy3VFpT8J6jt4x+O
ZsMQ+zdsdqCfsn3CrRucKAZjRLI+zdLEfiB3vbf/j3UKtLpru3/Jp6fHXKPPU628
Gx6q+LUlxGoDKDbdqipsDbcOEvwApALi+ObL1pMIXfQRvkWsvvpaWJEd3FCkwb1r
yXRv7E1Pho5IQo7bS98rCuejj/vs60sjb3pjH2gpHfa8PkkFcJ6koSvxQyCnmMge
jllfMI4tYBR+Y098nNHgXtuzea/A7JOVKl64+URiQJPtyN6X0YN1oHSUfEikCsSd
LamQCM3wQPrei/ft+TqW9Tr5Ov3maJOOQUa9HMNcJViNYr5SwQ1NzhZnDx+NgyEf
H0vzo2w/nqYvYCERuW8+poHLxPwQmZ22UFHpiSMWTbnW213okRsjisyQt6kDkcZU
MLDh5ydfpoVjKxoOP0rQfcnXc6llIVynH9q7U9YQg7U/oUFNKmkc2cFPsAE85fbv
9aBtoiEjB8Ou0K4+XJc+zaFyd0TnJ+iXlLBm1qS344IQfVO9EvrP4j+dpEMxDJAE
EpXMgHE+4L+1ocsKVbAyAANLCaqylTOpx3FVmhkwyYJTFLRI1EYKdKXLKJT72qx/
8xY8bh7RK1tx8qgMJaS9P+V88L+r/3WvStgZxgxZQFrMz0v1BOaPL+MHsZtOnjEI
FaTxeZ44e/h8sVYfrAWxUX22OJ/YH1fTbr3LJD3aEoRP7M2/tzaH+K54DGMSqGWb
v+kbH9NgVbqyPNXsYDRsmRQ7zbeZWp7bQWeEzZ+Kiu1S8glvvrcIimOzpQufCRq2
mYR8u8aoigtNetBRaVUHm4YJElicpSJ9Kcr2Hqa1a5VJT9uCNtMXW+1u+9QHvETN
EH3t9D+nfpglGXh2MRpoehPJts+NGcjSzxgm16DUrS3meoProPzC8QgYFJx8RmPV
zUBvgGVJ0Iz8idwnSSDmNx+v+W5rs1ZHnFMh3X46kPwaieo6xZbBP/WSHs8bb85V
eSBwRPkbQHk8vRjUjv7WYMBVWl6cCLFrUbB8ifuzXK+v59R/tZ7mQfbs0ULmTvlV
DANUkbcAsAWqAq4GlYwYPYfhFWia2AOaQuv9OhI0AwkZm5mBkVYrE2Lh4MchbZ4V
6ZsWDWaG5AZMqp8mlihAckxKgguCAj/VURRFOatUrXt2PGGqwAcejFoRJ4i2GWxC
RLml7j2GzfOSqUkojU+0sdYpn9o5yFP7im6aKE3bYqHOcflgFzVZikYlMSB5fNeI
XEC6dnYDSIDhEnl5PUUV9P/PP3MWmfdpgbNO+OEFrjbkDwyjkWQlgrPi6W/jZ4b2
rBbC0GpJfiHvLO6sHK1ZpnyMiEEebnLymwIxMaNnAeC6TT4aC/OmbX8HqbEL893a
f4bICz2fuNYj07GUwi4MqzxsWNbeuAf1RABtiqTY7ZOVJaH9hAR3rjJ5IxWA2Rlr
fPrBn9FaFeOQrwH9by9mqHb2O5J02Pz99Fn4l1rWdd0xWXtneRkpYov8gtZZMDTM
aT15MctdGTqh9sGNRzyGwkOzVMxPePzJX75tCybQ6PHI7Opoqu0VxRhfB0kEU73S
+uS7qFpbvaVeJRcMjlLEANApB+zp2nFHSjyZTB3W7dJT/CQ6dhxOd5D2XjELDcdn
/ZxglTzuURgx27foYj6fcWDMTG4MvIqDHk0WPllY5nREvDbJtJIUWqE3do4iFkdd
dbRBRoVv2S62SmZdh/woGwvXSzPiGmzRftzAq9kajK8sstTn32GkSGg9INlxmbn9
T+e9ebnbUCVeI24ff1DnUYqq04dy/c1egA6QQ2Lk0pEGFsD4Lzo7HUNBTwwpXPU3
XZM9VEJH/gXS7l4XNwAKDiEB2aBHzzfrwg6ausX+wabyKcp7Mfb9DQ+4cjKKa36F
mcBHhSOoP170B+ZeXwcv4BcTWHPI5gYA13zsjZQ8rbZn7khJWqq60uQugxsyJPp/
Ay+32UwtHkGsvuSSwVaSmTMKr6Jx7sFCTyjFvtnOjiit951GZjc4i4yeogQeDGGC
qkF5nccqK9ik9JyppIfBCXN4GMxtTm64fT4TwU5kM2HVdw8ynS0e8RLbGomE+I88
+iuNSoAIrf6eMQ3gigXK0LJ6XmboiJeN/K8u3lXNTLPxft5rtJiDDKUtJpNowphm
LcWU2vFGtI5/KHtz/R00I3LILDBM/KNk5AfMIboEMrW8t6MQGq3MP/SBtu/pHp39
J8ihMKhRDj9Eo2mRgEYkwrH1imzqTqR9PEwNrrL1OSyiMb23wbmu7Ljiz77SMoX+
QM2KR8GOyhnA47SOwoUPxXiPQ0QVCK+Sj6/1yMczfLNUPdCSkfklp3bm/6kTclAn
/5OQGt3zjXolvQbgRPdQ6wLDVezLrqufy8YSTwtV19Bn3l6BNrNomeUJEnNaOSra
lPqNoYTMj0N4s2srqK1KBU7qS+OmW88+YObJwE5t0X0PX5qRBOCGht782m30/pr8
t0vndIRqd4gXaWEREU/0pcaXkzZsvD2oI2E/EFL4vuZptQuJsU6/DxFkmYYU7dBY
W8mh1/QqDgJjTXBazk5LwwNViZWDUA1bbHlws92sPgrz/0myCcheFAkzIYbxzf4g
RibbYGyf6OlXovxKWfXCUEx+ppYTBpLBDqQ3qYngvdASOjcM98nb6t0p6Ap8cIVJ
55KqJty52UaBUev0F/QJ4+duVKyDXVcp3bAAG7bksBm+1HjlW+F7fN3XiyFfkT9q
t8qAn/QivlR+Xn1VPIDYbsyWQgoQB8h5aeBNZkYTOMkCQeRGawqJ0ctNYHm2kUcM
mDS9WJw0yMBoN1zWJ5yWybLFiIuLFzr7Xcbky2vzA+A3KDFTRcM3MyjA8I4DA+aF
laR7K5OMHe3AnL9HC6bOa54RNX9Ax2f3r1OsVhBTidRBIy4PO1yaIP5YYyO1aizO
osiPcD6tKqzm5tM80WaoLXHxGsL+k+oALV9J/aI842sgOLsUgmoMFqL0a0cgz6ht
MEbjguTqS2J75bvaITZt2FP8oT+PvldX0A5VQddrVpBTc+m844rJIBkMtsHV10fH
a9ZGtHGs0iZ7MVAsx2nLbHFbyEhyE/5OWxIajTRbN9rLXUW8HPkYXLMiDimzWAAn
hbYCasl51VKY51+5BeZfllFHX4M7ICBROdxhrsVcvlVRzz6lJBuRQJJ/+B5AaHN/
+YhjXH/UbOcWx+OhWthwsamGAaHZn1SjFhamZO3A5vOBhYy4w9c4yeJReA09GaEl
oPAYyk/Ex5XEZRLQdzS3aDVnG2M28xO24tbD94lAswl+MqHRQY/rHUvWgPYopHa4
rUVbMvd2jN9tSKczRiYhoDn6AJvMc1DhLLXsniP+u42/+nbJUSII8guVOXITIVkS
HR1KzF1WUTruKERFPiXpMGpsi2bZMa0kKzou5AdvIKRzVhzxe3JzvQV6pTF6gWoo
1ugqDpZS7pIvnCA0n+4PfPEHRAwIOGb+oUwXDfJaB9pb0YPLWBITP/wx30ta7O3k
R2YHilmHg+VdYPn6mhCQFIgiqH3o5te/olcIWmRsE6iQMeO1HMkJJDSj3+lu+LJg
o7VeGr69eIFsskRoTH4wQbGyD868T4wCXsep2250gdltcYpQGN3pqD81PnVOIcJS
dDKWV+vZLoMoQwHhji8TN60sloAfFzo00Uiv5v4rtojXFQPfvagay3hNPuYsRW2w
6HpeHHXnbiIC/sm3Xn/vrZcp6FBlWfeSZ1/n/qgezBsLIbpWNAOP6ukBHM1N1Lnd
pu10sFON3YZ9X7tDTEkMWBQjAcAgWbnDOvtg4qd4jocI5DOnARIyo3H3RCqiX6rq
wD85+4blFmRRj6zVq1BEaY0fkPkfBdiL35GJRGU21UDxd+vL1WxgdHvU+RSNFv4y
K2FtFcCPWnHlct5RgZr9K7FnTI1z2DsuAAg0WfhPhF5dSqf4EvKewbYpvnYVGDPM
XQc4p9BqRFT1ITLL1Jy8Z4AMO7LxZfxvdv0oewzwpgDWoQG/X6CkAe3vbdw7xgVp
cQHUD1wWkX5TpMYc/RxaWkNt4zJBjSpo+WDuf6eb9ZgJ8bgfKOojuQgDGooG6sBm
GuRJ97lqL05UBC1YTWzJkgpH9WU9rziwBACPB9h1zrTxmUE+hRuKndDp/wm/YakR
sOGRW4uAc7w/96VQS1FrjqqciNvsL+PwMOkrRVkIh73fOYCY/2sd3Pnd7sjGHhfN
UVI95F0xvOckY9UGHwgqVqFQdUfUK5jmHPpeXRL2VmSTdH0DDNozGTwsNkteBUt8
eSU4MvRhIqnK+SjjhJoRaax5p52xsNXIDBZQTUCi8fkbVm44ZRGX2GfAG2pGlnXO
oECKBftE6yjTwbApr8EUtQ8YPoWGFGp47GRAPCpyiiiDvRUoij2k6+SbS5U/yGXr
UwwfAaYXZjAc2u6NfaY+LyQJ5rwAt4sX0bOKsu81N3cftgh+0Vp9Cwq5J+K3/c/C
iWlOUmDuuI3hVOLTprXzHUYMhprIYLW5zZmXvlShXAoq/9XTlENbyWnYq+rzEG8o
cskslqW1csmqvtlqAwA1DBNNCe/eax74HZ7tvQpvpn79d/0Vu4VuoOrd4lEYz2Q7
io0EFsdkA+bRMS71o563f2f9dkk6OugQnXhHX0wT/7lUZbyI1YhYYtI7Bob847ms
4Qc9bAF1nH/UmhNArQeSM/s0AFHwuOHZY/plNcl3YwYjDJy0v/RqKiBE0UaYr7eM
ZBcBc2tbtBmy13nVjwzv6uWDrv5clhhyso6jryd2Giw0iNes6ea/IRxZQxJqfN0/
OJjO0+hiqEHIxckqeByBgC9dvx4eqrhePSSRFoiQyFOOlrhspD7mJj/HNa7GeXrB
FvXLFipxDnaPkHgiqmnhF7ZneROidMdwhLchiFqZqBMzPT6jZhBRQS7OPFy6L/dy
5dLPyuHs9h6cMRnbNom7Sg3RO8dEQNARtrlwyHW0Xw4S9HvZRZa8DdwNhhWQ8ivX
MEk1Jj5sSfcFuSUf/rhyhlC7ssfSG6N8Y+RaeuaclVuFuBCYG+xCCbKEByZS/ZAk
tFaB20PDavPvBkRYv3Dx5dEPLhw6Tv97nlkIXO6uJKGXwTDFtWhMD2//GVDL06Nz
SGs3B8fSCzzLQ4WxDVqq5rEbQ1kv/Vwh+aFk2ebHDC4vzdGrN8/VQQNMOzQUeW0C
IllGR4qH6v2w/OcJiGW4Wsnwmqr1shgavLrxh5G7HYIjHiYv8sfXhlDSMaZpBZA1
UsqGGTt3dbtUUqcF5kybYnA0ah8sTWfRuHU06zRvNrWMmlErATj1+FIpvFn92OKz
d3nZreFHYDjMj8Y1rMWJKZFyCouNT3KWF2DQBBOEviQAWcot6CG0vzuT74vNBTrp
ivJKoSdeaJtL2rWUz7YejipFcWPaclnKJR0GYdq/n4MFJp6DfXhN0DODq0w0+d6I
iL8z+xOtae+UKaMmjw4XkaLz8+bPHfqJtfKDTH7k0JCWHJKrpQE8FmMwPowrKBEx
hYaiITroL+bQ30LL7pKDV55i1uD2xzqORQog1RucwtYBTui6XFkkQm08o6eKfoAz
yHdqXNh+vnodjfswqRxl4CwkSmt5rcjIvt5cgKX/xAuKkIwBp72hn8i6OhEUMjGL
MeuvM2CA0ILqL5X7PyGujJGSMHLLqoZHdwdk8ugrYMkw1Glnux/KNV43tFipxY8g
sHrJ05Y4MzYFeFV1BhIxUZbw3nqpPj8zV8zz3QoFGfwypoUg2KXzhBvxDGcsU9Mj
VYMk0FiEylYEzNbtPEsXbm6dJUD/r4ZK4b9eEEWNiusy/pTMdDpc4i2BaM7584ce
e5WcBbapLhZQQSvzp5cUY/r7yhniwxsCmZw5q431T7gPV78ko8SMai5C7xOg1acK
9QLOlpkg4VkWAjCnfkni1DOMoXNTnZWe6WTlCKJN6wR4Bn+MfvYdfG4gOzPpFKrr
Ou11Qysb+iw6de1cU44u3Jv6F0IbIpIxfOxVm0l8zow+d086ySJ9zj2GjCrGTB93
wgRAWi4xP4yb6W1aJnz8T0oc4YsNcEnMVvwUq/pmaeQ276NGxzInCUq0C8Vv8eMm
qrGMiDfRWYS97Bd5K9tF5575dlS1wokg5MUNcQ+U/mbOK3bu325JCQoykqqyPud1
DZ5DyB3lH7FCFdHqJrv/fH0PThU6I3xUdQn3+o0a1m64vUPgVhSx0rlop2PmAfPs
VC1YDk7sMhyWbCYCUpSTwZKUBWs9ccr1B1Fpv4JtjrAp2gM2MdzomKezSLijZx0S
/dnK3nW/HdGrqDIr/W/8wD4/bLYed1LduUQrQZyooh0zzZA6CNrWC7VFYd0DbnUc
+Xpb0zgc0w4R8se7yshBtaFTp3Cef780KCknS/0c/NBKarH9VeFWGmuIVwI1c9zo
WikMUi/YsYgh++ZZ2AsLozvU+oVy5pLQlmRXr2hvk0P2uWecx245DSnS3jjRRLMh
XIchZRUXQQ0IzWo7+Hv5fJ4QwUNjaz430N3l+bg5sHPAZRBLBioFmIf6fkUik9Ds
Rrxiex33FiuyUzdWDzKzFDsS0VG72cxqlFmPUY3dos4kU+ylX9rnPzAsHHx/TP8t
R9dGKoampEBO5nfCsH3no8oMbSnOe+yeWlQKlhF3XV3eXO45eowYANn3IREIiugA
xMAFoBz4h9loMUPttTKM8/iegPu5CONIcYZNHcoTX1639vAHqTWlKqPemIYD2T8e
QLB97+9HvuHKP+9UflKAkYe93AjHQul8AWN2tQ9PjDUcVE6wZiKaLljZnhxnhrUL
OiygorFxaM8taRZkOiRk0glcP37I9Uv7P1It+3aVzyTda9moLmtrHd8XcxtcnUcw
jUFY4+NpSX/dMCv+3lez2DAOY6OIHLyIOmRMiVC+QbecCo5CbrdRlZuoPEFsSM48
a81Z4ZigUzKjT53xbPuBtmElo2J5LHBAHLqf7O04kTL3d0niWgIJ9J/hnQpeUOiD
2P3b5Y3u1lYlgEBInzDpnFFTXCUyEdHmp7YghGA/p8GUy8sLO70N79+thRyyhAeI
ZeeznnjRMmONguvUlmcyHlx2echtG46U6aCPh+liiK6mlq16m8kom1ZGr+Ed5N8N
c4I7+auf3ypgS2kK0lCGLjnNnI/Ff5L4AYTE1MJSuM1i/RxVCpzeFMudH6INHXK1
uz8ubi4N2jJpkOJiZDGfzTxGI6kzKiV5TH/qJT3S+ZBkcvAJ0bGzcaS8lc3pWHmJ
NAsgNmZ3ZrDeCzIr5sAoyNMSg8AQYG6hGgnvJ59Q9L5Lx0dez4L5iHYMw0pJeZsp
cV9yjriWi3Yu9qlBw1FIs+XCo0HYvLRqhCUyPcq3Ks2z5yNfmupQQkpx14FQ9dUT
2RB9GP/XpwbJ480/DRG5Fe7g2JEb5IdvSb+skyJYiYsvdHz/kIlkplzll0w/pePc
o33kXcWNnqKV0aBWrPe05TiSYDrDBWwihYI9xAb8Q3ER2CakmTadhp9TM7u42AoQ
KAz8JCDRpDo9jgJs4w4mOktb56y+3/PL06QaOOwvrjnqGCszyTJSHKYpFTnntp1G
kHeg6vaqXhIBR3R2fkaKCVPkDqGN+BXys5jaLVdUnHKtnV1ISqEjr3ToTaI/28LU
ghkmutpbVx7ZjLDWMI0BmompCdhLsrSYtPxGNIpVgPHbXavGBV04Od1MNIODUC+k
PPozldx0gZksq20U7MtVx1a4jPeWHGlGEwBwSv43WvuyPcuTm+YpuGdtMXl12wb6
hUye4GqvcpiWnBHL54LBKESXOSNUWUSPuOxWfRLvL8LjTC4EffYSMPIF7sm12qml
4H0jD5TgmKyAAPtNf1nuShIDfqnELSrvHWZJZe/29ift89V4mQfVGfpgDpDJep3H
UEdbx04qaD6BRw5pn2tiUwYQpJXcOGB7isprycgctPGk4zNb4/BMXl0NiF6TXi5a
e+0wosYfhTbFM71ga90SFVwdJ19Nqfl55gY7/4WjrRjK8KDF+aC3qcB2tRWsx19z
6Z3qB5vaQpOC/vcARJEIlPBLI0Sfytapky8jMfoZT8sBmkpcQzPmnzpZIbbWd3Wt
0wlqIfS61ufneEEofW2q9Il7eMp0m5Q6VraxqIV1zUa3ggJh8eNV9d/YxeEQLyeK
gPJIWg0IUif7k6H1/vqQ+1105AJ4isS8PtNwefI36wiLgD+hCeBHy0n438vDlvfi
malukP96NglPojraBPm4xc+rcy9WCyezjHWfQGaoB3y61G2BkeSw/GvpDX/YS4d7
TtowBLWIB6qTbQU0gT4s2fJhR851stRF8z4VbXEFFf/YcElbiiVBChOf+vvB/Qhh
3M0WcF/pyzI7PnFQxQZvuXSX5Sh9RSnh6g6A+Gl8L0IJ78sAuZ2Ru2XgjkEUBAEU
/gRoFgnnxoe/i0UEDLAB7cb+sJryiVSswadEowtjI+LxZTv0JZ27pHgNjIRs8OCm
+CKJxFuRB80amildU62IbzDKwDUj99wWEiK9OmGbbqbjaMwQ9YCEiZLWeH0Gt0Qs
GCDO+H6QxoHsXxNtd/n/RWJ55Z25zjzNCG7Vxqyr05lKEy1GAEWI6CW5a3m4hILU
8WOM+FDghkiKMroQS3aAmYDDRnI7192VeAPSng2BsxDcltQCVt1C9xQByMgeTEoy
gb12s3MVgt2fEz9qyAOswCqSOJz9qI+tBFjyWJKiYnEiGwdrSEJjY7lE6Kx1IR29
wpQGQBGeW5ggaHTHSgpq7afTCd4b07d9iex0vziNuK1N73UXDpWQc503QVO2L+yz
UabVMwgQm8B2pvZITbh5KLZ8lTQiZ8Tq5R7Y1YXWvezW0IsGdaopGf3OXZvuWZvP
N+PcZOoTyiXY5COwTvRtBda++knVpxZNBL9TE7HazJ1bt7Qt8iadcs+VQYfQSTgf
XRHVZ5Ie9xHA5Rz6u4jZb05Dg7TgYTgFXVOkt4d8zu4GR/uUXpwUJINZ14U/YbI7
sOKC56dL3mjzhWxyPbjI0XKPrK4OOoMsoyRZTwDZiI9lwV8XKsLEbkIyeX8uVy2l
xQPbrC1JzHjYFII+OqA98uD61Ey2tzIclXLPiy5dG05J2xHB+qdz+jjf2jL1TTv1
llqqwcxIxB1ReW2N7//y8T++2Gnz6FViMXl+TK3AEAiTdU7J3eVtO2revCMhD3RE
JlgFlXsG4kxE6LApT7Nqo5xy5qQRXPMnGNA8R9BqOV+nB9/4mq5af6pfWlfiiVd3
6oXavsvfkCIB/FAhklOWVPolvixxpEU65YZ4rz/S3S8jlxAsAUOnac8NOhq6vl1O
2xk/88MxMXfwY6mYAgjgr05Yyn2Y27lDrkQllTSPpFk0l+Jr8TcnVi7N8qc5sdvD
yKRtm47iQOQpugw3rbZcxis2LhIPGJ3TU6xf+xEajlFBI7z5ZNXR/KC62pfWccZ7
tzOVU70ny7vnTHoUX8PM0avd61f5rBkTr1y91Su9j7l81mSzb69vAujej1akEPON
m2sGcY30aJ9baP5K+H1p6mS1/z2oLouCKLoEnDEDyQEYX4+2EuSR/tLmzw/nS9bE
XZCQgBNOIbIoUm8Q8WlqXJJtjZECuesvsnGJGFUUvxGdS+unI1pZaXD5Zz6s583g
aHclST6KpDS7JqKkGwmetKNL/aLme69nqaYtUU5AYm9K3cfwYnZpT7ZCZ/bzDcwH
QWWgLyedzNWyqiwmFX1/a6NhYBmBAQ3hyKYI1ahIfHFkwEGs40axhjh6bJg2LujE
X2r6CD74zzRrzChXHO2Bmnm8F3wRMwtfJnwooDvPDKpAZ6ktp0PQjXlBlyQXXib7
XWju7QrS13szAjmjzhQ+QiB+BLR7yVyO1Z92rudIQJnix1mTj0ZkudJ2+Zlv5Ire
mg1VSlRY6VGYTwL/Keh+igYRLv9JAbQm4+uKDSFYZwL5syTegigDGSN0mcgvnNP9
CWYcA0bM2AHrel7EvNYbvgwQb+QNQwqJx7LwcBn0D3gudrKq8wNLoPBRQfLkaeQ6
FhnqQM2OnJ6TdFeyAQnY4H72fHpEf6xYoFlp8IUdRKIce480/l4PIq3WdQ6dNY9t
EkruTK711juG5jTX9oOxERMAegLykfkXX7Mqbeio6aJuAmU+aQxnrHRxp1vNKEeC
44wPRmcQqcA/0klKCN/UYef6t+FfmZnhbOmZA4CmrW0qs0HiNn+DD7ATpHf89Frx
mJeZ5BePrGhZfqyZulPksLPr8jWog9XS4RPtxYCbIQ3p/QzoyX7y2bLuE/moyrno
hW2kbSFhXapIUWNolMLQyN0K1ozStidbkBU1QiwWsv2zTktZRwt4crNS0+jd/bnW
ykp9btsAtNxZ6/fLXY2N2DPFr0vvM/Lj4WaCymBxkrYF0w9a3PbK1T9xmkGp7iQ+
Nxo78keHrO96+6cHTbSolGLHJ2YCwq/svpElEfjUknj6CVDYr70yzKE/OUrb3EtW
6YjKCDQ5SFhkcRZaDscc+8TPja27Ya+EZ+XL5mU2TXtiDVUSEI0N1y060BQmW2Yx
3DF8LYIpxDAlwi8vvuXoxehSFvpsNkBRnI06zQ0ane4q5NcBHfOagcCr9+fJyPKB
qaglBXWs526IxFtEIEAg7FtQoWJ22s9s0/O6CUag0GOEpulyrS4E5Mrkq171m0Vm
/q/wfz/lo+m8pQSwzu/HH+2qbwoyogjPvvZmLE/6aNNzFa4oJtRLKiVZSuFuF3iM
N/YG3vXKrZdO0npqrFXfTENne/0wKVJBfDSh+lyyt/4t0EuY1mVK8EcbqdVQsPZC
mEx6SapNmqJUwbDCoeF42Lw0liUsyGFoI0l5b7B849RrK0XANVRECVU5w333c11C
zvk5lZH56erqyHCTUej49rd/bZ7f58uA/0e2lKdAp7FUzzI6QdhHF5ycUHZOyEQ1
ihPOxH48AgjCT1RjZacs+1Ueu2P3ahN/MKfRjUZrhmTxkNtrMOahBOMfeZwHQkNy
9mu8i7ERwUHiKBvbS85qe1+kg3HkryUPNzQFJ5aBc1epqtGRSeSGqr2c4FEuy7D3
Zutf+0r5zf0l7Sv0wPcGmdSQaWQ2Xe+uZQKPqbidzBU2EgSFssRPfsn5EfLqFSz1
S7iV8Tnm03yLVtf9riAeLj8/86+X6gBzq3Llfn7K2MpeMl5udUlKmNdujGHifxIO
e6MHTEAXRgh8sRRAGjQfD9Gpa7Hokny/bo5xqgVkwuBqck3LUr0Q1MRfJ0smD7rw
VpT8I+3LEbcDauFH+MjzNhTGKq3KFd1B3gs8fB/maIZCRTgkQHxSHCA8+YeiW1Hj
R5UNxy9sWk+5q9xRBwDjODhZwFqBteYmv/WwLZulb1T/7boPk01RRejJlXIeCXGG
1eI2gXA+KdrPK1gz+Fw4VItJnGKq+7SVC0OiaTWjYAuvhEzBpQLn8lm/xk5lqRWi
84yFeYGodCNxciuWbQMO+5d7LHKvkRKCqKfb0qi3vDheIYFtQiYiRzC6ml7fHJY6
N7Pm+Ad1coKxy4Gb9mv3j7agSxr9+yTSf8AAJYax9oaE90PJJvEO/+iww2GwZrOn
991r3wYZemVrm/oBxQ7bqZz9dntx4e/DO/Wkb7JKIC4wJcMUUGHlqID3f7hwEyBd
q5Ect3vvG4sk7JhTOuxYSJcT9fVATjgrjpW8iNHxCdGp+QcTJsBIOIb+RqExghx5
ZrH5nJbtKjEut7aD2AP4/ei30CH8JhWUabCh5vNY8LGQp44ePnvXc75eEDPaWPvD
+Cou/5Dfogw36nQQeN/7S68/Ex2xdGd73SJ7D12aNv9lBaxq+G5ZSwIX/2HJF7YQ
/mEsUPP93UfC/zySGRL2PCNw/n8Fasr9EGFjXuA0b6MtMBsBBy2PP8nJkAIxnY3R
gL4x4B+SdjnXGAnBBT1be/Xo5SctoTosnT4ol8gLqUrncejV6OcDQ9FCy/o6jOH9
5mQjvIngG9CiWsXHGMPqUssr4xbRxwV3mSasAKnOlB7q52NeTOTQ8ZUf0QuoRK2J
TPgU0/NI7M9AjVdaq3arnh7MvpUpSNVSOFCKH2TKyWZm49BjN+vYPW/8isgj8HHo
DyvnP4gk2IdI4E1sf5MXsnCuZXLnxwA8/AxDLNp9Jj7Klm1ES08ATPe4WfsvzK0G
umQH17GHBMQAr3Mt/i9uILCvixGIXX83k9oPi1nBrNTl6Q06tLmViRnwR0UU+X5h
AQcrEDUx5Mvk9RFaRRqTLyGaKxBCqQVgS+bEPXJDJGqgacXp9KeAeesBxGn/oxhg
KhrgiYmT+6wkaqQjjWiAylKO5YayXnwQVR2oBznFsKUlIlZZMCOgXoBMRP6eXSt+
dTjQMLSb7axo38w0vGFPhDwftZ8IrfRq0B2X32CBWWslm4wVZLkJCeWQeh5pqZTj
n//H9jweVrHOdQZX95yYJvx/mX6ymGQomy3DMt8nj6pfZma1AAuydbSHuncGCZvg
6rapgBRAKlgGO6pbsM6pYYeQ+SQxD3iQApYWu3J8TZdcJnM60jlhNu+1pbhQoOm1
UjMRU/EyovoTxDw4XWnLdVHJ91Xpr6fNAeGyWSBPm5trX44xN7EIw2+M3aB2c1DK
ATnwyBfTKaVZBC2kKWbp6nNOHsEIHRctmU++iSCP+ULlmqYp73kVdeD5r02lbxrP
xPkCMQRx05+NBxNpNVGDHhDafiJiui08GmVylhjWf+bOqcb9DwPGqjZPAi3Hx1Cx
VjqqSKCO2vEIGIvkbwTphHjdbC0HSG4IRK/FgTeS+DAevYEf+++EAE00D2Y1I/cT
JsQD4eLw0RjHKT093cgoiSjJVWnYtFJAY0X2JDyx13oerGh9t7GetMfZ3ATwX7Jc
43dpd297aqR3LsIpQ5/ST18hhfPDsDnBYunu0CURh3ZjEXQAHNPYgHGc3xMo1tJ/
H+kMa0gkntPR9ibRRDC0A68tFpP5u5195/J4yumpZYyVyEuyFIixou8AVt2ADC6l
nLk7y4ZSCDrHRyh9Cn5auTt81o1Q07iWKOwY0IM5dVHfnp6ZVSCvdLyYq8qq7TqS
yhh4cLAGqUzclxYtVRmfKoLyybdIMPXNLm0DSFSJ9Td6FPdx20ZuZqcElmTFXACc
a1Y/Duc8XA7drWh3gRowtCKuF9JquEwfkJSuLd46lAP0pGWs1lMQ+Wp8nnc+29PP
eqNhW4DrzNJNGLbx5uAJECzrwKxkkACOlmp07Dt38Yj+UREjdf8UgRI1UhxvJ788
mljfmoiKfDlTlrKqRTPpvy48AqwK8GgY5eJyJC3qKEYZKc04OuRS1B8e6F3A8yXq
Y4Nfsffgo367CcIZLjBbBiMtl+5XQeqDnfE9BdN4hxigCE0a89wo0mNMkalPBjHL
Y+nSeBXu2gZLkxiSMZGl7001GQVNTydZTvCuJpmVbuWzquGdw5TscbBxeK2ikxOM
+69gQwlljn3tJ2dD9w1PjlHTUedbSYKHBOGwE8eHbT2EIy3m8MqzL7GixumxNjB4
eyMEm802GNFkwtA4BC7MAzxE29o60ePpmgva7abFDRk/hl2/tpcXgScPU6ynretC
gbUsUpmDCHMs6Hk8AHCfr4SF1BDze9KlZaGwkwbfcqtLr+jowfxAkxhvzMnQp0lz
hOCnyhihEqk8CX0vIQS9eDIETnuz/NpljaTIFgm1svSD43O6Cgg0vh+rNuP5gzGB
6f2+YrlKg0lybZ2RN14I9oz25SHBbM+eMEMOAGidZWAyxYKWeVCeajA5FTK5+nVK
2yicNqPB51Vuw9P3av/eXIMlFBSRFPslP/kaWUSzS8o0alJlmgbWvlSw92yVQmfr
kXhGjxyQF1yQ5V0mIe1HdBDENfcdzBunmPHLE+4KxA0WQk3P29PwHqXzBylB9mV0
IO2AGGlSK2RBnDYXwoLyNOzQ9SzYUYRV74ljB7ZSb46c263jxuT+vnK0R3XgnB4s
l9iBFRhJ6hMPSXdA4X9D76gALLgZqNobfbqSaJ+y9HufaS0fpYQVgdFCx43In53f
oAN7au3cIrhb6VORlqmDB6bmkqN/j6roC3CSaRKvshvqzMys3GL1JIK3t66J9D85
Qv66dLH15whcw8TuT+LA2FHOrULieUNOLLaBvCRO8MX+KqGesdjMQwlN2JmeXi4o
2yCiDUbsKaqo7M72Ynj8jvPApo5g9myEffhG7RekslLi0prMb3I/ETDB5/qzClI1
ui5qyfmQn7BJdzB9ckZA2X2eQ7KD6g+GYR1QY2CbunLoLo/8QUFuuxCysDiClNMK
0LR0LozrzuOkvniiq8jOSbjHu6/r5VlvICzrdi2ZXYYTpZkna6k1nDBIsxQGxEbD
Kuv1fgown8s9f69lm140jUkMv3HfOl6tMTECpaQHtYurTASSYjVMJUiY9xx0Uy+O
Lol+SI0/KND67wV5+G/IyJ8mdoU2iCdRz17eZ6SXmeCMPbSIFNCbj+NRzYG3AB0L
X+14z/rSVeaHnBKu+cTWwHtzamUhdsnAfEZ5FOm1SIURA3Kw+l1zBmOAy7lLQTpe
6UtZjTvbcS7D/m0svzLRZjTue+IGVlQKcCoEIa8Q6PFbJgnUkqXxKOWOEvV7DOlU
D7/88JqpDqgU0a9DHFGRYBGdkZExRgElUGm4VZr3Sj6UKmehEyNXifP8Y7LBlBAS
+fk44vDb89e4vBAWeNabM16R+H7XVp14/GnttgqnV0fmRhb0fS6Zs2nHwjsrC3eF
wcAi8jUT7rXe+il/tqXGR+IuNo075vGMamVeeNhbgoPJncGjnyu1d+9A/se6/XzV
CMkYhFb1wTip/m2xOtUSfV5dTNq6wECnk0KKeetBWOvgxIU+EFWCBQ84gsDaag8f
KJD2bwyIyAFgD1xhzORXjHTOtfeFC1FMY6137Fr15E+lwqTj2pBy/YF3Mj4RkJWh
whjVdHrI1eFSBMSS2YYc0X+mJbWE/R87PvcH+oCsC7jZbqD+nlZu4iubfTf1v9P4
RJb9AMvXDZvsTdCEfDIf18tPFiPm+xKyArmrU3Gmjgx3X9iSGN30dnetaIx0PxD3
gGvzv4S3RFgjBTaB8NEv389bUIxHOrf08Tv6nE6VhLttkTKHjwtbYqQAyv1tUKc8
7LudM/HvUWm9e+kc4lByFRm/li3sOSytk1SNUEmpinMa9WdfZybF1DDdMCpDKale
oTO01HwuvWAyEviDu6h2lFPwVE4gy6uWravdafz6AG2WmPcmpSQqjgk7DG4CQT49
J0oHUfraZUn+uX9FxWps6CC0mb8k13LqL72U5EDR83qgDjTpbFoOFzUQS97Y3Rpr
zeurU+C7uRWmDJsDfHYxiebuTDZqFa51aRhpXgADSKkjh9JoXN3IUBIGJyV4pR3d
uKzp11zXEZbwrX//woUnJMW5xgC57O5bvKwKlsv2vkVyPVbVz+V+azwbSoCKywox
4VrDSsh+xm/8CQmBcIxr6bR5i68QndjAMtaP0V0YLYczc8GK1CakzkzuAGuMd/Aw
q0RQLeqP3tk4k3SbPyb05ho0jzxvzDOUAVz9TkQZTAeLWfHajGWVW+xkZNqabEAS
8UvJRstZ+qVzHxjcC66gZF4tO7E6AiTinWpW8CW0EVEwjNUerRrE1mjnU9sTGXY/
1aoO+WBeFS4Gp0nkYrcOl/MwMmAZmx5N6v1PhsCRa9amZSrJCenaGE+ySTdPo9rn
/RNO1rFzi8xiE2s6ZFAUHS2HKGsLC6ky1cdsDt/cjwr267uA5pM3eNSx6sAZkFMn
cMConOSHaIAyLnMUSuUjs9tZ7vph9/Iu7nGBMpbWeAWA1m8aTOpIXHfbt5LFUzzL
dZImA/bMmpFo8d+LUtnC2/VP8KjGRTMfGvgA0mmpJ4NRwHIwFcilvckV3JflwCT/
ZIa9e+NEuZ4mNSw6D6LLE8A8y6h6G/xd11SW9Fb9EQD9Q338PCf2ILt9HN0M3VAo
Sqf1TZLGCOWROtSBaJF2YtLwhHyv7AV4bLz0WCIrHX+rOQwIpbbB3VvOOCTkkXu8
f1NabOu1n6vEdPucgrHnGtjX4vkdexFeJFPZ4rLwMf4TZOa8IY91z56nv3ADung8
Jtc8a3vkeRmoMlOqmjFHiZgATJ4qDw1S62xMTYRZvTllbOs5N7Y91Evf6NiPTNn6
o28wJELL+i7/yo2EorebWq067pEh9IkMmYqDCHQsQ9VuH3DKOBPX8HNlrC9g3FZr
sN5tFKw7OB6Bk5ChLJA8I8dz5bTJwIQPKbeoVrSIIphkygPy9mhiuPxVNvA/hvRo
l+kUriMTV2qtxsaU9b0a4JWnMHXwMWXFZ7rodZs2kFFAfNsFiCf1DKzcpAvLyW+1
ii5SPKg2d30N8nKIurRxXrDh/nCWuQ/XPGWpVtumZ3IVTlXt9jAdK2XAKKQ0CpnU
sydV/m7AEQ2gRC1BWRoHep8H4k+TMptTODA7tPcgPtIYlESxS1MlmEG9JooSi6ro
qlxSJnihpBlRQdcZSRHMKqyhm9aq/2sbMENsRGCIdUh5Sa+2KsMIxd1eRNeLQmup
OhcBYbmM9jmolHMEBi4rcqT0Kv0YlCE63PZL50FP3DsaoNaBmC33M7KQ6wXQw95L
BlYwNcp51pi4fM0eo1bMVseaelyg3wQbLLZqUtsqeRq4QHtIxQYtyF0+2dRsJAl2
LOgnxjgILgNo6bx5Vdxl3f+RY4AIqepc/05VZzVkaFpIXUpFiUs31zUDxKVYIy8f
jXPn1rL1rYrJrDk+ScjP0Bqi4F4yORur/x8Dq5Q9jmv9pv+jIdTuFHSvoF9OB0gc
XaCfYP14gm8VKa3/1XSDV7dJc+ZcjlT/WgIo5z5SHcfkY1IANgKdckjhkcBtPbv4
oi33E2TqkeyCiw3ZQkCqvdNQgRZSiMgbulrtuLIhDbB0h16iNr0YQBRS0ped/zJa
CVfNWnAuAmVOpNDJKQeo5bHl6sqGK6NbIYsbPWCpYrz5kMlaQuFMgmM6qe2MgCLS
YxOgbA/AF6QDY6fqzaFb3fL6IcglndRyM6boATx4tHaOsiEy+j0i5Ios3BAsxjIh
MvxR6BLNZRfsiWMXFQcZR+zed4N424lgTkUpJffYbvm5zfqWaBq5FFGxP9aUif6P
38DTIrNqujUWmL7UNMp6HOfYK4dR39L1xvef9ctwGZwK0PEds1n1GVKYzOSb8S9/
lWxrKsZ7+5q1OEwBQHkajidpdxA5roVxqI1kCSeqssmcuE1SIV6BXg2bY1nhjBbi
ODes/pd/h4lnl3xj4VUViR+CBNuEbGw4iT+5/gryIgxVcSeNpZwpMIcqtw3Zl3Dz
zGWRrzreQAV1xA4apdGcBjTztWl3x5OjTT8F9fvgh4ozeglixN3L/dMuNckrcJs+
MWVzpNv1saH5U1C70roj5r9Se5Ym9GUCGdKDvxfdy2fsIIth2imijvwdm9mcLGbI
zcWFBKbtYZ/pjcu/6BQNif+2TGy3Fwp9fxk/ozfeG4LAoAvN67Fze5hjCCs8IYPp
qpL3vNDGk3Iv53jPySxcHZVJXU0NYvisk8faLBhdx5igHadtsB8RD9S8XcDc8Bza
HnIH7eFg/DN1oN25s/YFXGNIsnCZnofkLFWkd2E7Pm1JA/Tw4SErm3FwYfEsA4og
MEcvvw//DO8y04t1Z/EsSMIv41KfZsrZ8TwE6VuF764ARA3k4QF9awAbFQfWxG6U
3H/OXX920Y6tOK5UIy3V4kbVy5/QbS2SOpTPts8/VlSxMt9HCZwZT+Gk/BmtZVNW
nNNnls2gBRf/scYUdoBZEJQg2Cm6kAWZRYagRnR941G39ZEeouL5LCV52mYGTVsO
YaMntpE/DjI9wdEjbe9ddXQu2JgQzwY92RGaGTaBuyidt7q813+BeMgaSyqW4PR3
Xzhi1k7UXlruAAqWb2rEdUHtw6i3dvn4yFI8X69Hj2n3OCJV8A8eAJTQg6T+sQFh
bEkjg3yUymHGx4GiTx2HDXlnqC7i9VSIUC4vEFTyULNbTeICiKAeLYurM0bzNo1v
nVtzAkF5yceebDSB/L2/5eEukTfh2O2409e/ElgBa4PP0DbauQYvgRUFrt6O0DJD
kMe65YDKB53ITcTEHyzaJQDgYLaNvGxdghle+z2zxuNhkNTmeQIBscUl8n5sQtS2
yOzLOZTuxB/B8lWI3CZD8cg9fRGRuIXj+zOZkzPI2dfmTZg+00vIgVGxuFlLH7eX
QSaOmEhJbfwQTo5ZiMiEijiMbWPjL7fTaCnSsZeoV9Bb6oLppTjqnomHoc3wHa2G
rBjbXzMTLDoG5g0TGuLgMdxqJiUSSHog+V7jmL5k3PXltE3R0Gsbp71SEYz0xMTr
`pragma protect end_protected
